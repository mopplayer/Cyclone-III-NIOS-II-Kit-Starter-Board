��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_�����yn9��r{�{i�:nS��x`����7�4���ۜ(Jd59����G�B�I���*�m+���F2z���>�;��u�_��̿�Z�f�|=*�b�7��`f�J(�|�~׬�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P��Ms�¦.e�	EP)��5������p�nJ�8;QB7���f`��ə��	���F�c@~�X���߂M�U ���[vƽ֍,X��h�\��	��������,�}B��F�� �|�(�c�s���%���C|S�[��͸��|~g��ڪ���޿�aܞ4C)4nT��!!�'���z�o fu�����^���g�m���2��a�Vu���d8#� �!����e���V�9q�e�NF];��Ր��2��P��z�p9��vx��2���#�b�:������HO����t���Gm������3u�ݲʭ�+�緺�5ZK��E)�����2��E�0ʦ<֧��9LS�Or�KM}�1j%��en�R�b�z��s�A.��m�xp����nÇin�`<p�&-8X�Bg�Ne�(�|E��T�&� rg���6qn�X��X�L�b��g��6Ŭ=)�3�I�C\��]9�.n�4l'k�`�	��������4�;������{r|_Nn�w�<U��=&˔�9� Gcp���ь�;��Gv�{�ޥ'�+�B��?���iZ,2����z�Eu6�����C�hL�R:�z������;nBs�D�}��8��w���j��2��"~Q����y}%���i�ًi�`���_��2��,[QZ��O�9D��8|_�c[��b �X��r܎6<��s�E�P�V|������M{�~3�^�\|;f�@[��0͗���!$�Q�%W�z3Ň\��pu��i[�/:K�����Q�w	
�6{4�:m�%%�,�?��7�4�P;	d�
���'�E���=��Dy��|2k�.ז���Q,�^r���<T%˯��;"��)�=�������V�!��NMe��e��6и���VLst�nX�gӞ���� �㺂o9ݯ����Ժ.o�w�a}Pm����C�pD;��Ƀl��[���ws�5d�}�u���o+�T��3��UTlp�Z��F��,eg
ނe8 �!=��l���r�Ƞ\V��?�S�2x������v�m��!#�5�aA\?"kv�Z~���x��Y�x��9�mLe���O���/z�t�?�>��_7�N�wa ���Q�Z���@�S�'|6ba��<��tڂ��>�a������{�V<7h��-7�c���{<4V�	?7�����P˶O1X}+��q@�ZY����=���u��6��!��,A9A佒�s6#e��ܴ��UJR�h��)�5ÈV��Nu=�oz皝��������.�8��5~�H�6�[��2Åf���w`h{����
�����ulA�HWצЖ��ˎ��x|=3Ty�-��!),�#я8����(��R,7ALzޕ��ڝ���ŀ%�W�d����-���K�X�֨�էss3��"7?�ȑ(c�jQ��џ�x��)h��T�� }]�Cr���Z���E�2)o����df*r��`�^pS>�NR������mM�"M�0f^��Y�S�_�d�]ڗ���b�c%DȠy�A����	�v��^e��3=���V������J�zϏP0�g��V�-Ps�E@u��="�%Yۍ(��˃U�>7y���vM
z���O!�����dI�@�De�/B�S�Xpw,҆��0���udKͦwM�
-Ӣ]�Ax�LL�����@g����E��ʞ�tq�5��������y���*ï(��?p�3�h����ӫ��֏񠞟8N�6)�yN� ���he�1��ɷ#��sn9J�&^ِ/e��F)�TQ����~S�D�N�$�u9�S�؏j�0��������맨p��((��N��M�ʣg~3:��֕H�g�ޱ��� ���%BWЛ`�f����#*���[Q~X��%��>���(KݻPKg��KM _�L
}��NM�J}fƺ��։�\[�>0B���F"~=�`���È8P�zt{� �Ic.��=;�62�z'�Â��|�e)<?��⟩�Jh�$�rl��"7-V��X��>,���`��B�+��E];�֬�+_h��W��+�Ƃb�����X�M����(�j���"p�H&M$r2r
$��~5�  ���:$!:�=a˲���x.~���/�ZW�ߨ^TLHS+�z1ZeC�2`�J��*G�-��H�{�7{�D,[���0R����p��Ki�2n�*���x0�%z��	]2;�D�4F�칣�N��K=L���� \ג��T[�8�Sa�9�A*�j�^K,�<՝�Kjx}���	�)�	=�y)̷vSr����.A�#�;E�����L���5x�ph�f#�ة�������]�!L-\���6,��z�����\;��3�/���#)WDT0r�\�G��"�����i�v��/dv/�3;{T��?��+򛬞�Π߹��q������C��48:��V�% t�>���<kF�c9�m���8�to��P�t����Q��+�=�޾����V���Kc�#.�*[`�~@�z�����l���>@���e�r���O�ި�N�c߱9�~�Z�+�S��;�6� z�������w�{ ��_Hs�fNiU���w�z��̴�Ga`��˯�{IJ�n޴\��4���<.�C
1���Zr)`�+�9�h�OBq���*���Z�8s��gvl�0*�"$a�v(�Ȳ}�Aߦ�ű��d
�m*q���5Ԕ,�gy��BS)�Z7 b<V���??�W.ZR�V�s�?�ﾫ�-�eWI,���0�V_�(=&�n���/X�8h]��C�Q2-�﷏�k��2����"��v��]BR�������5��a���g�~%���37��Ћfͨ"$�n��4�P�l� *3�9-����x��"���7�1���m/�A �A@�/-�Yw��eDyl�t˫x>YHp_1��A<ʲQ�K�*���[��]�/�>�ә6�;C��6F�]0�N8��L
�1�Kg�Y،w��S�;��V����U�"��
FȆL�B�����؏'�b�1^��K$
��yܯ��|qvq�tϖ��s��
Uya�>� 40?��ޡ�y]RU�q����i�&6��v��<I���p�G?�$��wj;B��O���8�x*����� �*B�[�P�#?R�b9�o���JT� ���yq�|��T�n:�s����m�ߌ�/���bs��*�ߖ�d/�����j)R�Ѧ-J�}�� �J�>�*��H�4�},��lN�A��_��R��S�|V�G V *���J�8��>Q����Ȃ�%N8I�ǻʉ-����fe+`*�Ǡ@Su�M��t���8ך&`���Ͱ�~h`�+�Xe{��ƍ�����N�wQ<���T��1��!��"��cqE��]�$`PJ&���:�A(�,k���َ����YD�Y��Ht��֒�pq���	���7� �Y[�nݧ���#��v�4r��&�r�]�+Y�t4�ĩ?��*X���Xŝ��Q)�%�{\Lo|�"�-WȚ.����ڄ�
G[3:�\|�5��n��
9���!<��b23�������*��<*��ZS���պ�}�I�?o�Z�!�����[S<��XƜ6%j�0�t�8��[���]���:V�1��a��x��� j��A$�̈�Ib>�TW��/�!z���D�x,d79���~�[�����w�I�_mcr���1F�/쫻>�z�Tﮓ���*tz�&���`$Q�7%}��`O�sF�]���p3�h��x�j��y�J�����*�u�z�s�mO���QuQ)e�vp�r)m���Ѝn��>�L�T��90�_�Ă�Y��VR�f��k�a��Rɤ�U�t���v;��Qy�@م����o,����6,���� SI̘�t�>�Bg�(�"��@�JIA���Ͱ�e�)���;��K~�ˁ���{<Q��=�*�a���{
�v��&U���|GxX��U��E���cMAhB��e�Be�s��]B��	�\� �H �]ٹ�EQ ��d���^�ژ�2o���s��@K����0�9�gs7�>bN�T&�G�gǹ<�$rIw\C��L��{�7T�X���E��`o���Z���ݰ�֞�m�ৄD�E�O�mn�6jЋrE��pS�xbW|a�Y�H(���.g�_D���0��2�ag]XBz,��h �����0��p��=�����������.^��h5�Bէ�j����]�8�l*��q�u ��r������=�t��gl��2|kߊ�d����;*�S/��2x��?WAvcPU&Q{?�TS*��U�B|����<�1	(0�U��%�e1e6kg?ܲ��
:Qf��1�LQ���s���-�1.�?�9az�{OCհo��=H�B=�ए�Ųc\�(��#ڕN���j��3��yI��Q`ҜX҉#�������6;�N�%�եmU��YoD6*���Po�Y�6��5�,�R-`gfQeK�KCCdg��]� ��D���{�߇@�k8y��c,�`$���'�Oh鸋%l�K�4K@ϻ�a͕YG�����! ���9�����"���ډ4v��9r�"��Y~��z,W�oT�ͷ��]���֍ͽ�׵'��2<L�('G�b�H"��^gg�c���n��}�C{w�&���\��-۝��}Eӣ�p�k���n���3�=�t!����?�����t��ɍE�W-K��sc���V$�C�X�*�k���޸�د8l���K��[��ۙY�:/�B�ke���Sm����9�6$���ؒ�Ճ.}z@�8��T�8�Q�O���H,��D��Op�2��%�D3Ӯ`p�K�q�&a-h�}#^my��k@��<��S��&����w�c�\Kkt���r�+����1��6�fo�_NKF��^�1�\1�x� �v�)���`���1O H��-�zyQ�F�&���CDؙjC9���v��AR��}
���x��A_'<|�׸����Y3T���>�:Pu�*�;�,��&�,���iq��d�i�׍k��B�D8FY c��3�����5�nPi_�Ӽ��aJ0!�A��l8%�}� M*�ϯ��v��=w�a��ڀe��X,��Yբֲ�R�?q+��]r�ox\�$p��V�+����m��߭���{Mh�����E P�K��*��#4y�����)�T����&i��ۺlt��/���
�"?|���C����t)�f�X����~tk��m��-i��&��Iۯ�a#[��Jd1m�A�N��/ 	;̃�gX"��u�D���^^D]ކ	v��Cx+��׫����ǹ��\,e�	�0���[*��G�6JZ۽�QK\씭��<�d�mp1����p�a�>d<���q+Iy��q�Z�0�>u]n{��1�����6l�2�`ti<J�p����N��4e�WE8ǖ��_����A2�*H�`����Տ"7��S�O첻L��y�o�ܱ����,�UsB8c�=�%<���b�RSә��q�0�J�&
Jy������>���tg��[�s�6	 ����k/���>�J�m����-�A�����xe�Q�Ô�G���C]LЋ�K�0�;T4����4�dTU��Zϗ"�c2�����邰�:d�O�m$��FF���$2�zl'�U��[οx����b���4��ʺ�6�Y� diup��>'��[��R�nZ�ȥj�V����2�Ĩ���hd��A�7��c,���Y/>�gk�L��)XC�5n�����a����A\eUsj�-$GX ����n�m��!���܈�-��x?7�����M�=���4���ՐqeZV�I�E�M�\�/��-{A�8:�^e�ܸl�$G��e�+i��cL�\���վ�j�`_�H�S���,�!����m�8�dg�8�p.�A�d�n�䯌kk&2L��i�Q	d��6�?V;��Vq�4;��2�!���oB��5$DX۔N��9M��B{K8a�|��%�B��]�%ïZ$�Q�{Ms�����c�z��a0nMp�p %h<��Y`N��SOJDZH�o�x�	$��C��>j�n�����{}Ր��o��\�eW	�M�6�#�"⎺@M����`��e	Ҕ�$X2�p�m��]�!;N�5�p����V~�Q�J����_�h^>��N6m�(��/6�=mS�1��fZ/!K�z�p8b�*���Ѻ.`��
��y&KS;�asSj��w�:�*�qpF���]ǐN����z[�o��i�閠z�9N�aYx�khpy�p��Z3��Q���w�#^l�b�-C.�Jf��o���vX�ᆇ�;�����������ü��@��^*�#$(��_5�<��	˱�����;H����'��Y���ણj�xa��g��N�������X���b�'<S}B$,���C~DÉ߆Z��E1Ro=8F�6`�"�\
�Dao���gR��	I\r�j88�k�ɍ�!�Ƹ��M7A��+���)�4VjT�����-_��B�|gn��77(X�=J���|'��F��9�ڝ��x����[�r�'��?I��Ύ�T��7�e%�N*#��C�D���Kl�'�x	.�C�v�y҂G�^N_��#;Q���͗������۷n���ki@�SI�58�ǒ�!;p�#�hM�4�:�ϏE�OH�Hx��t�hcޒL�C7�:y�2��a���%X�F����OB1���#��~��:u��H{���^>�����h�=�	@���T����� �nWy�!�ӚS����[j��A&��$WĢo77bi���~���ΔuGש��D���zM�n矸g)V�G�b���`)Q2M�u���M�_N�p����o�e~Ŧ<��������MNpH�u�8�uE��p *{rB��w���
S��S�|[�0��q�/��~cp7ͪP�c~�u>Gc*h�����6�u�AV�4�Ш�מi�(9�,�M_��X�3�5��Z)�Y�8w��0mZ��݉?�v�^q�0�������/:��r%k�)��W3Dr6��//�^6Z�}#��^;���K��/�C/kC��EL��.�+n�!8�j��؎4i��Ƙ$�#���O�q�~:��-aP'6su�Ak�^!�D��"ҹyv�b����d�����c��\R����X���oj�Ɇ�@RzT{%����`�����b����D�:s�u��٭`�˽�vgE
/K:ͅ���a_-��zS��p�|�.,j�1/�;���\��$�-��`�% �d�}F��ۤhE��/�̃:��N)��o�}��,{� �����¥�����Y3�u�
w�CcO�:f]Y8�A`h�{7��'�q��'p[PP5��)�IB~�	��ʗ��/±�p)7SX��5�CS�E����!��>�IEt�;O->�{߂Ʊ�Li��M���kc��Udi������ҐW�5L1��-�qP?F�`�V�R�V���-�
��!��Z ^��kū�`�8�N
�Ç��[Ǐ�g�E��9�����hª)��K�x�^DW�}{G=i ~*/��gXS�{6���0�u�oJU��3�[:4 4{�kH�2u���_g��PK������F�=�ї�v�0��QB��s?���N��\l8�$~��TD�������� %T��#�����*Il�)`��Ń�H��U�����j 4j��1�OD�f�uR�ˋ�&�v1>�I�<��UP�U���m�VJ��~c�"k��ڕN�p�X��񶖳�#I%4�G\V:�R��u���\��$j��g�-D��7v%�b�	�{)����L���I�����i6D� ���ЊGm؄�־��^��@��c�c��D'��7�+��ݛ֨G�䂎���<1_�=�]-�~�(�XȦ�as����ZY��ҽh��Pj��w/���g:�m%ƲBW�	�G����,�5*���YP{���	du��_D	���s�pvI��Py���y�i'k�9M� ���uè�@�.m7�<4��-�5R�p�
�p5�}80=�5Ƴk����Y���]� #o�>�����\�z;(n��7+�	�}}���b�X���X` E�������w�-6I;��zG�E�2E���O`!�yޜ���F�|���<ixt�4���*���R�w��z��)�Gྟ۠;M���B�l���"M~S��2
���M}���'\l])si�?_��ߨ�]���[��C�D�eB,3�$H�9&Q&h��_6e�},S�f$m�I %��vO*\IX�� P(����I݇�O'�\Τ�:���lIq�;��V^�_�)뷦Lé>kH4~?�KC���6����2VD����*��f�p�7��d��?Z�½�d�}���Hl�| ֪�gZ��l��+1F|z����ˎ9��l�
�AC�&����W��B����ܲ�$U�(a�ϫ'�?�wA�VN兪v+�*�>5�un ��$�w�ϭEէz`�0X�C~?#P�}. �ƼԲֺ���m�/�>2������v�͆ gx��`�9s��lRYn3�G��s'�����l�Ni#kY������h�l�PP�gT�M�Zթ�f˫��LJ�+Z��X	������"/���{����W��o��?Й�;+�4|N�c����@^�܂����v���
,M9�,u������6�v�{����9��9 �pnUl��8��+[JSԕ!$�cW	�]�}�u`CL�0Oq�9b�c��Ҷ�Vu���}�2&̿m�v�J�~���Y��ΕңG�s�z����9����Y�1S�Mk���
�!�p�4��>����)�e�`(�B��~؁-�ճ��4�5z4~P�����Q��i�t����g�G���
���h(��h�r;B�i���+7� ����l�!��ɖ��� "Egy��;G3/
���4�`�����Ph��o�Z�p�CF'�u[Y`wA��M���9�����	�-�yf��u�m#|�Q꬗�V���ǙY�l�Ҕ��p�"}�NC���?�t���yc���CP��U~�#Κ;�|Wj>�5<�)�ȡ~ ����ޡ���Y��E�%���y���'�&l'Ek�/��L�L�<��JOMM��:��~y|�>��<P7�޴T�f��[�"��Y����Ӣ�����[�E��Q"��(/��Z�g7Gx8+g1������n��xwT��Q�}X�S�aA(UC��A,D$��DCt'�X��{�ǂ_�axq>u}Jo��b^7s&��H�����v˧Xa�ՑV{v�I���̩Kj�����w��Q�O��9��f�F�7�!T�օj��zN.m�}�{j�%��F2c�56�C�д�@�:ڍ�Y�;b���d�1����ۂ�[��vW�縃��;� ��,uI��"�����3��M�N�k�@�p��lZi�5jgp(�k�%��#8���6+����1p��l+U���a��=��Z(��B2��vt:G��M����}�
C4s^�����D8Fu
ST�K���_;Ie\�����w��X�^d�� ?O �Yq9&��2�_�~6&@������oL�
�����N�[� ����/��)8o�C^db�)�&��'����F�h:.9�VN�w` hHQ`,����n|�I��]�)^�S�r[�#O�^�FS�(r4���	4	��b�F�q��M\��Z���_'
-{�S�;@��:��x�"e����3Gɼ	�R#��(*i�\6ZӜe%�r�!&�1�����`��_���n��g�-5NO �!݊!�>_N�=pyn%�Сl�',D��UL��2꛵圍�Q�xN�n��9Z��v2"u�NƮz��գg�cEzQ�I�+iR�O�"�D��-M�TV��Y��r��r�n8y�*��O��IU  �W�4dZ��h��K��-�U�/�h,��� <�����9�rY'u�Ң-.�O�x�!H�؝�Mw6�1����V�[O���Лb5���)X��y*:�������ʃy�������*W�K+K@����tR� ��g�����B'�}II�9�M�i �vD����X_��k��B6��Ыۋ�Eo_k��?��u��]����;;��=�y��<T��el�v'�W)���i,@]Y�������=��RK���{>�����/��,��ZB�2����𔆻頲�@<Ǽ��Y��ax/��C���W��6U$�������|��U�#�[/e@1�j:��L��̝���JW�"�}%��Po�CQXO�?�J�ӗS[�ä��GK��q�ߴ&J��_)]` �万q4	�գA"�։ј>b^���X�sJ�q�F�<}�}���l�hm�e9;��~�v�u��p��Z|U��Y�n	�/���qd����N@���ʦ��l�K�\K�s�논��S}9 �-�B�;���rxD2�"Ty��42�x$�S'�"t��dd��&�)gPG
/u�NR��'
	��ر���9,1�E���-�0�X����8c�#IZ�@�.0��PQ�o�7%�c�fl`oX���Y^�pi�"`d�jS�?��){����Lh8p	�u��ouN��?RI&�+��¿��؉jR������f��O�9��������$䭡��dT��b��Z��f�M[Cf����7Ӭ�2�:��i��`|��#.t@Oc���!��aĔYAȿ�uլ�T�֭*z�^K���t#�汌p�3ڵ� �Ȃ�|w���թ���&�?g){B"҇i�TN���=(�%}F�S���z8���{�����E�Z}ove��B���'���B�m�:�(0y�}\ z#��J�/�!O��h��0�$Ko����;u�tBTw]U�Y���T���z�<1��q*���� �a�K��wلA��
�(���֣i5ɗ��E�m[bN���^�4�J�I�Ͱ����=XDG���劻�%`h�o)mlH��V��Gc#`�8)"��t���ﳹ�x.Z���;��\��h'���Tu��q��Jњ�Ϝkb��]c��Lņ��K���Y�ؠߋܬ��� &��cZ<l��T��%���^W	���]i�?Q$��95����D�)����f���0���l�	���NA;��:��3ׅ���b`��!�HڨD���� X����m�Մ��w�4�]s _�'�i�$�S�k>5�WF�"ފ�'bp�:�3�΄CΚ�N[S9X޵G�yT��2L_�\��W�q��{z/�x�3P�����߱���f�.����䚑����b���p��$�e�Q y���ti���J��d΄�-t-`�n����Wuj{��ƭ(R�Qrd; X�\��J���2+v���9D���K�3
h�i�U�CUײ�9�h >�E����G0�u�˰S�$DlX< <׫Z�h�� �����x����.��H���Dn*�����7�G,"�5�t����s�뒍�EP鏨�S��z$�5�.�_�
r0����U�zP�r�+c��<XnL�������k��OC�BL2���p�AQ���`,B�72W�w)�Ca��)��^{0��HD�~�v�r|-���TQֱ�@ALd�@�]F�_Y"M�^��N�š4��E���0����)�H��X����̚#��Tm2�t8Neۭ0o�l�J��_[e( )z��5��i�4�'!��������z�~�Tņ�e����U1NC�OG�*4k�YB{/Y�\z���칔q���ٍ䘰ॉ�~�X��6,���HL8�tx��"�ߓ�����keAzgWy���WK�wx���^{P�4�k��0֕o�[{�@���@��c�oU���._fq�4C��"��S%���j ���&��F����UaW��뜇t�EP���+�'WI����^�`��v�<P��O��)�I�6 �틸�Ƶ�<;�^�|��r�n&ǖ�_ ��z)=C��9�I�c�o�t+D[��g�H��Լ��7Z
��./�Sd�x�s�K�_Q������ j�y�]	UA��?�z�Z��n���V_��+V�}��l{���9�� ���X�z���\�6~U,���/c��#��ߖT�{�ʽ�Ds ��fz%iL�w�_]��;l�c���k��_�Nē�P:v��N﨣�.qH�f�E(�mS\�X]('n��$e���h62=�C���"�%���]ɤW�9�nJ���T[	��-�[�����qQ�s�D�������p4m�C��̙��^�1τ	;dSy��f����8|���܈#��X,�_��:6��gs��(�z~�Sdl0M:��9�����Y��C	D3�%|a0�r�e����u�Tt\�7ʲ�ũ��0�	gz���@�,����\,H�+�X�ˉh}�j�&q}�00!���̔�GK�9r|&�+�i�M�2�M���!10�P����~a�ff���
o��˷����"l��W����~�����'u a*)���
L����±/cōG��O���uxR�1���VuO�՘iN���~���Mt�a�!�� bʏ����@-���M�<�u�z��.� tt���
s��
�0����~����������X��Ś�B�#ɣ�f#��� }�Z�1\ WD+��G �6d���'�J7_�B��p���V�≛��(��e��G,!
{��+�*��X:7d]��ɭD�"i��A����r��;��o�3��'q\��%�� z�V�*���p����(&����ō{�vĞS��{IQX3|F2����A4����@b�~g��WZj��K�����9��Y�"�E�KSe�PO���3DߤV�כ�%(�K���8�kITm���(��j�ݳ�rS9jE�47n��~�~t'�6q@c�~J&-��S����na,�� p�f<=B�ɓmO&���R�E"H��iΆ3׏���/.�Nr��I����ݫ"&{�>��K@����ƒH��M2��b>g~��lJ$����ڶ�"p�U��y	(�ԥ�W']��b�	ڲ��%IlX�� �l-ަ�lbS�u�1}���X�:X��~����k�|W+.x�zD1�����Ҳ�{�����-x�����V	����Qgk"�sp�c���)��	,�����v�*"�06�������X�C�q%���M��zy�C!�cЇ�'l��!)F�k�x\�L�09pg���?�MH;���J/@ԬNƯNu�"5��3�^ԅ�ڏ�k��wHG�TIm�V~`��ǖ��d�&�(�Bk�)��@�=����Уz3�!0'�Y��?E�ʹ�Jn>�� B�"�� ��je�;a����$54������Q�������$=�2r8J���jo�:� ������sg��/��5W���[��[_G7u���Z��g8������������u"9kj��*ؑ�����a��,�� P�W�D��1$� ȋp����SԪ�L#�d��^E��Y��x��}6�;s}��;-�,��+3%}ڍ�Ɇ\GXs��:��w�ܱ�̴�D6�NJ��Z�!�G�5���i� �ʅ���Ey�E����Vu��M��w;������X,O�n
p=�����U��)��J^�6�@������ �ݦ��u�9�ΚKߟu2�Y�e;j���_�ݿ���r�#<M�)�`[�\��2��obZ����'�v���s7�_>��jyw~n�`�D�c��/<����x���Uٕ���Mr����eٳ� ���S�u�L֮�Mx�v��fB����4=ډ�p�B[i^~�֛��G?�w\��w��ot��҅B���F�
a��c�ס}/u�U��/��D�V�7��0�85�G�f�d\Y_K�z����0�in�>��.Uҧ�F�sXB�$���3t��'���!8�A�5� 0�U�$a˿�bV�-}I�ol�N�0<SKq},���D�߃7B���-��}����U���G�x�%9({�]��dzm�;�+_4;��p���U�{"ƭ�-ZKGs�&�O�f�j�5w��`�s*����
?�>~���j ��~�1Ϳ��x9��u�xD{��4>�P���Hz�4���l�eY4�����:�#�1�[����%�������F�,bPE0f�vxH��ꎪ�O|$����U�Ν��]�
����Yο��Jĝp�ҭp��Aъ"Vh���j�� I�m>%;�<͈n��ͦ�ʨ�:h�Qe	����@i��8d�[�Rl�%Z;�	 �v͐G��Έ_+.��Þ�ͼ�U*M��6�N��{���&�0�W2
x�.t�I����p{Hw2��G�`��պ]���8d�r�p�3¹�Εq�����3�b�Y,Lw�S������r�{JO��g˃��v+>@�$��H����M(�g����(
C���"KcgK�6�S��hH�!
��o�x_x�YSѐ4<e����o�͞nF8��c�%t�-+|����Vk���_�TnM@������ك��#��cf�,������B+}���U <�H��0=$&\��?�f�n7ioUD�kES�t����~:��U޵�����3�,�# n������">�|�ē���e�A�[E��M ��mط�y�ey4���4���[�r��{�,(����5�T�����U놩m_kIi�`�Ѩ�[���P�� G ~<n|����o��MK� �2&��;��u0?Ɛ�9���@����	'_��|�&�|�q-/i
���{J"�b� ��Ci��-gf��N���w��N&�໷�G��]�IϹs���FТv/ȣrP���#7����MAGfA��"酒�)�		Uk3W���^	���٭���~�.��RE- ��+M�᷌�t@��9ԛLT-�LB�@�O*�}��G����D����3	��������&E�e�����4֐∿�� ��aYr����w� rQ�:�B����A\;�-��=�WZA.8��y԰@b�J�]?���=m�F��c�g�65���gA��v���.����<~ ��ఠ�p<�ψ��s��ku���ih�����{mE0�h���Mߊ���o`��.�>�-i������	��i}�T2Z;GQ�9��4
F�|�I��K%GYF@�{�&g��7#3�mS��P��S'|�_�ւ�n���+�|9���2�J:XZ���-@n�9@`�]�q�F��yf�pR�����e�ϼ�(����O�S�iw#�L毕������5�|�������%h�W2�o� ���͟��8O���䩰[�:��w��*.�?7�>.����\˼~�R؆��,�&󣐷�\��� (v)c��S�*#D��~�r��c�m}JC��Y��YE�B=�@oz�&s
"�Tf����[ެ�'�m?�g�5*s���|�2
]uQ)wv���0O�O���绪��r����q�(@�7� �՚�z��wi��6�q���P�m�:Dp��i�)/1*} �c�s��93�/��1=����=��_�M�#�%��Ϊ�7�f�"Kc�k��>�O퀞}�fx��� ��Hɵ��ɑ(m�dM�-�X W�� ��k��	.��By���W��v!�����t�?����5�6"�	��Lqۀ�l{:us\�;�X�R92a�}��8z�?MF_\WK����x��^o��^~vԔ��m�_E,�d�o˙��D:��>��o��_��x�(Y�œ��թt��-x�N��"�v�?bs�MO��_{z����"q�%�Q��&���]r[�ғe}?? �{Z�2t�p]6��t�{��G���K�C��w3%җ�#ƅ4b�������u�n9k�-�3�%�#�b���%d9�_���Cɂ���\�+1m�a�=^�u��J�F���l��6���#��(����Piq;˅ct�AA8v����3�h�R&��]0ƛ���O��(9�(�M�n9��Z� ��Q��.E_���1�C�]�J���f�9���O^uZܷŲws)>�^\w���ʪbs�zFY�[�#��K�t1L	��W��	f�_�"T)��m���^蟈˖<� �uW�����U3�x������ީ�
u��C]��r��/gxE/�L0��#K�b�����3k2��I���I|�~��]�����W߀m["	�R�1��/2���ZiؔYWm�~�B�rF|��1c�#a��Y���~�W����X�١�e39��G།�5����YՉ�.X	����
��)i�8�.���ّbL9`8R�7�%��63�������N�~RԞ�"V%X��Ěj��@��ށ��tPPf}vT���)���%K�%���r�O���{����:�I�>��
�f&ϲW���ހ�$�@�CbqQq9q�$�V~kGL4ɢ���P!��_��x� '`D�D��1���62pF�8R��V��g��{v<�gPNb8��iW�ka�c
E��`��y���s�0#�/�s��#!#�]u�V���.M9��2o��r(;
�?H7M��w�F-�u>8䴗ú��c��%�=���HU��QI�#�+&Y�Y9eL ��ĉ��:���~EN��� ֻ�!wn˾&1�2�m~U�֮�S�n ��1�K��™ L�J9oR�@��p�K��V���az��غ��欻��������o_(�:)N�ވ��D�
�{_�(��w�t��I�[u�c������#(�8����h���l�������٢}L�֠S ܻ$s��=��g\5�".�d{Z���Y��jRU�?'���S����{!��j���:^K�H�>wdײ�`�'5�aY��L���gLѭ|L����@r�I+P����FYr&뵍ʜɓ�y� u�ÿQ�
V5X:��s?ɛ�qէN�����9j;��f�����XrT����=�
�q�7�N��s�.H����q���?`r��C�«�E6�9��pB���_]A��S4�r��\
?₇�M���؍��ca���.��;�my���S7\��ؘ�	2�䈞Ҙ �X�͵���z]���Θ�ĕ()[�_�̀f=U�&�ʧ������ģG�W��A/xbA����9�AƵ^-;��!��|�oi(Q��.�� *�Z�1p&���P��L�㻰��fP�i��lÜ�e�(�8K�,]R��{'=מ��,o�[ڏB�Q��!�i�qꇐ,����*��$\y�~Ea�zRp�g$N�$U�	�JJ��9(���s�����1s�A0�XFE��-~pM���]$�P*>���,�#���T���Eo5�$��'�>��4�u��M���'$BphW4㍙\f�ޔ���-���q���'[=������{PˍO2+��u��&Y�޼$̍d������XAN��>�n��u��ڻ�t�j�~��
����#B���6��׊ʇ�=�r���;
�D2�d�?ʗ�)�ʨ��9�A)�'uF����:c��Ũ1��OOR9��V,�?�d./����fp�I䚟]��g��F�#��@�0�"[2����;J�^PmV�kY�?��mwH�J�ɚ1���R����~��{W�eV�K�o���w�.R��kw2��7�s�v�>ɏ]�B^�r�I�Yz"��E0��ZC!Ct��<�}W�V6I��9���O`��]��|�v�b�����bW,��@ֱ�P0��={��Z�����U��ڎrZһ��%��2�|�T��2�j�D���N*;�	O���S��)�yk�5�ɺ�Y�?�w>��хX┷�Bӻ�P�MaW'U��J��k�d��_R8R對H���YKs�H�Ж�4�J)AɄ�e�D��GS�Q"�1�S������g�����������`�6r��$yuQʶH���t��&�6��M�a�򇁔"�0]���C����d��4[�VW�n��l2���d[��ɷ<"���[���oR_/�?�~�|��5�|�2��߭�*<�k��lg��G���G�5��稙�kё�AVw�1Ap���<V���m�|��4�T2�˹�BZ~$��i����:.O��ӯ��{F{_���Bg����x��패Z�3$Q"�yI�,K!�*�4t*\�������Z��'N�<�2;7Ͷ޶�^�A�ˊvG��\[7�/򜅳�pM}�X���ʄ〇�`����s�r�\�oR:p�ĸ�]Iy��*L���L���A�t��d���y�{�):�P
����v] ��/��$M�:�̻y�� }���BE̙�u��H���P�aA�q�P;�:�=�R ��7m�k�a򟟬�%h��d���CȆ���
V��$���f�����ѱ���Ç�
f��ˠ��ф5q�E�%�ڬـ�}N�k?ϼOo�u�W�83��_�'� �!ÌR�<��OA�J\Qj>��Y��'�U���"hO`Y3��>�R�:T�0U�jZ__��A"0�A��b�=��X0�朗p�����u��Ss�Ӿ?����i��c-�z�=��(���+�YoMin����crnn�Q-ekӧ�hk�M�(� ��V�Ekg��%�V8�ɵ'M� !�7+���`"Li����\��h��qJQ[Y�>粉�N��)mS��
�)�Ł�qi�Y�[��a���		�1�{�w�uhOG���S�_ΠH�L��������E3�gɢ�K/	���b�b�������g�a�m�@-2�<��n�ަ�nw��LN�Km����n8c8o����2ha����I'��v�{�I:����:�a&�B�l/��R?J�7���dn)h�m����e�#�����������x���9���5�E�nbe���F�c�|9O������F����Q�}v��p�7V�\�]��?-=5MG
\iu׬���K!ma؞����� -Y/��$G���c���@�G�-�YnV�maF���I9�f�B��N]�ÎU�q_X�p8�_~��@C/uv���NF�(�������o�e쬲J�8>h%:��X�o�bt�m d��(�^T
kJ����āL�5>�ʗ��~5���۵}J��.-� B'A�3�V�#��(xGNNQ��"B�h��99��.��nf��q��������4�l��޹����X�ïM���񻒋$=.o��S�	��TP�?"͉���>#�g����������t���p�@����-��S'�˔����\�_�m*�:ce�Ё�۴�@�M��L�,E}&����3�|��"-sI$���ޢ�е)�;�PPt������dC�҆�*N����U~��j��m&�$8�ui���Ms��r�3�
�u:j���ť�[�tj
1�D��N_��F��-#2,35���#<���o�#{|uh�}�EE�����Xld�*͓�ߞ[���[�ƽ,�p8#z��Zk��g���m�nq΀f6����m��]9�����uE��|,��������4�\]��ʾt�xS|N��/�����Bg�쐳��*:�AҀ�%���f�8���2ՠ�7)%�)5��ڧR,2�q�+>tKx)������P�h����<�8\��W
.9��2��B��i֔W���IV�孋��൒!*���4?i.sK�t� m�	$�F��E�q�<E��S�議��O_�G� -�Lפ�pO��ʴ��[�SŢ�e-������ӪWV�ew��T�OS��+���1�3\�;/s���z�W+
�|�*C�d�:1Z��w��
+��m��и��/�?)��z,�A����AZ]e ]Y:�ߜ�:�W�lx��~�"��"�y�3¬A4`޲����&��/c��G�~Q�h$b|��4w�eKSM_0�Tv�ob�]|�BXܲ���xd�|���p�f�$�"d��el`�$���3�����BkD.B�?<�D !#��?�������>������[ӮI��l��P6�,U�q��9�H �O��������?�&Dd ��4N�0h �BQ�r�G��v�k��� B�\1Nj�,#��Z��a�]���w]�_m��*-erw��S��P�ZR�z,��:`�~�ބ�\�A8t���	y��]�a�J==m�I��1.����9�Mv�]�'��x���z���@Hy�����S��'�YuS5�Wq�z�[T=Z#�>�!t���{�0U������E"m_���r�䝷��Dp������/��{3�>J�j����'�(s��#��A����	�#�>�f���/'ɥ�t��nd4ɛ�jt��$�b9%�|�eA@i�SE�즽an�v��U�)��㷎��1�G\4ɛiF��A�Qό�����o)<,:��Yҹ'D�Q��-7s좙0V�I$��.f�
Rh�8�9�*�(�􈅘�p������XaO�/Y8�
�0��`�"ȗ�_G\?{%K��;�t-<���N`H�_Qc>vn�T�;�U%�7���B�6����r����&J%�]~ټu�ŀ��n���k��*+�E���!��&I�
�莁�e�k������(.��%��jl�[�\E�Y����������TQ�^T(�<^B��HW�o/�¢c�iL��r�ΏÐ����T��牬	
}N��M�]i�r7����m�>�}|�~Q7��Rʐ]��s�M�U/g����g���0Z2<X&��+���\���㼜�	L\ܷ�w0�!�Qp���R�߳�s?�bW�N<������:��}��XUJ��5��3���f�D�e=��3u1"Jg���S]�7�z���8n2<-)��R�OE�Q���*%��Պ���j�s=02��l�V�.�� ��|�B�%�/^ �卶�zNa�N#΍'}V������?�>�\p=(/?��#�ˈ�B.{L|�U���󣶷�/��)�{}�B讓 ���U)	�N�\8	������s���\�g����j�*����$�W��c6_���F�"m�&uN���?�X���9�BofSF;�s�9� ��>������[^�y��y�7/U�Z	?���X#�2���~���{N!P�J��NnTs��w�oI�L�`^}l#�d^���@T��5O"�k�U^]ԤUTv���C]~0=0��i>H'-��,;y�@OB:�8�Yfe[����5Y{�� ����M���g�$����<C"�3�2�p�_��a���~,P�]�%�5�\B-Lo*	�n�J�j!(���e!�}43��DY��!l��d����Mt�\�1���Xk���h���m��Z���_1�Y?���J5�+����1�K���Q́�P�&R^����C���QxWo�O�p�٪_�2E��=��*}A%�|�QV�M��
�݂g%�(�S(�ǭ馭YC�7�E�v�^�v�ȉ�T<�� U j�V�^��n^..�����:�G�R�7`�V!��U�U�V�Nz�hO�*g�=�'9C@;Y-፝?���M'��Jj�D�m k �cz�#-",� �>)�.<��J�����"����wΨj������Xp]9h�7a�H��٪�ؑ]�\?7%�H"7�g���+� �bW���'t��Bj!9Dc4-~$�Yf�S��NHlD�ާ�i�bɾ�!��u%�=[���C�Á��Ao��5�(�:�t��7�#AG`�X� �b��:�:�4��x��-�3QB��)��]8%F�*�<��/�Ws{���#��k���I)��5~�H�������r�2��$R���%��$�)�
�h����y��M��H�r�EvH���?\�౔�7r���샢Ʃ���g�?�a־"�����r_4�N�k��:���Z3�-������t�l�F�PJ+�u��ԅ��CS �=�ڡ���TF���� l��EV��_`�d䡛�����W��H��Ḓż#�%�P����`�'[WO�m��>tSK�p(։*L��ho��D����(b^�Δz2��ƈS�'���]}�����zg:�ͭz(%�{�\a&�c�p�[(sC����
��'�L���-�$�wGX�Ņ�E�DEJm�5��>M��oٙ��2�����1�_N5�<aQ�H�@Ur�d��eLW&��gC� ٤Q�B�v1�ud,�e9���y�dӰ���όw�-=�����&������\;cE��e0L�(GOI���l�e� jX��ӟx�o���$��v�џ����7��[���]�򶇷A�]<��+s�:��O��Y�'�*S�s���.����'�-��bg)�i\��'�:2v��}2x�ox]!A)ӊ�h��@�rR��X�����JئڈcA�qF��;v~1�:�K��+�顒�N�0�W��X$�":����ƀ�����X(�f֮�s?0n^?�j'Y���d<��G�����h�KUٳ��D��\�݋g�����`"?�S
ϒїT��������g����l��;>zuz�J�Nb"'��b�Ί�T�e�,b�J�Xs�_s ��2�'��@��u�����Z�c���;�Ҁ ,���YM�9�1rB):�e��.hs����F_�^���Sf|y���e�𖧛�e;��wZ�.�͎/�ȯ�|i�72�R4�M����l�R[fz��1�.��vO +΀��u\J�zI��BY�Uk���!��/�L��H������U_x4�L����ɗެ�!'_�J��;�v"�4���C�KW�r������t���}ҍ�%�:����5�j�>�U���?���$DI~�B)��v�� ����[�+cx�p��馀�F�3�W��µŉ����R��5HrQ=��p��2'��$�X��M!� ���%ч�T��8�oV�Or���Q�s_do��9JA��U�W�;Ei��ـu
�b"�mz��J��&�Ӎ��ҧF'Ы���Ʌ�6�I��qȭ9G�ʋ.!AJ��Gs� @��:oɫ�dYB<�3pl��'��+'���/���ў7Mb!���gl�X#rD�<'����a�J�*�i�*L�NKF���<b0��n�v�wf�����I�
'Au/{��5�F;�m��ە����G i�ġ���L�h(�-���N3�� ig�Tf:2ȷ�U����00��@��J���C<D��iE�S��9�*e:���Z^`����y/f�ˌ�]�K����ԯCb��?���V�n�Q�]��g���M���`l��N��V��y|J��h3��g�O�Ck��5�M����m:m
PėꜜS�Ke�odkXS����$�ڝ�=�W���s8J�Q�ͭ�3�7~D��WC�>��4���{��bi��4�0���y�������*P)��,�O�O"p��E�H2aRb��,��+c�,>VY=7�4-�3{�0�,���$f`Rz�j�&���(�|��J��w��e�VG�\t?E������T�(KLF�^���5���׫��^�\[�k9]�T$Mx���;m�S,W��jA��@��~���*�
b���@Po���[Țf�AG�wב��b� �c����$��.][�H_qx��:���1Z=QDq%}=��rkrҎ��;�e��~PT���D��2d]~^}Âq�*��w�*�d'�	 �ZRO���_L� �ܥm\��;��C�~��`�����l��}Z�wW�5CwX�^)�*Æ�3;5�r���NK�
 �o�ԕF�PST�2��b�ꛡ��!p������2�*e,N���H�GC�&��*�}/Zk���c,v���+�h��4��]K�e/����wJ�{�ɟ5��m�!Z�(����J����\G�)�ЖWU��F�+�H�>�˸m��9�%�t��U�u\|�[]��vDT�v(����}�U&d�A˹���1�x�ڤ7��SJ�ΌFXd�����$TU�oBx�
��`��˜�2W�[�R�1"��R�Y�=�	�Qћ;^��ip�� .�p��VnK�~���+j��8�MW�|�!jj�!�*s��m9j	;ز��K���R!�d��ӹ����U&u=�5�J^o�'���Ukh2�m2o�}qq�&�^��|�C�"��O�T�c8���d��{LM��t�LR�Ľb� ��%���N���÷�t� �^a�v���tS���yG������\3���RH
[�f�8�ΛP����S�X��S8Ip�l�0���)`n%��ڭ������Dw�:Z�rAd��W�&��%lC9�O'ˠ��� ���S�Cd+�c�%��R��z�b��],��|�)�8�y�1�hF}\������E���)Q8=tީ`��<�*f��K��U�D�]��?��&���/�T��B~���b%�+��ڮ��տ��
�%�-��1IJ�Ý�*�4�Ú�S{�K���.���F��b��HO�:���'�&�[\N�.7�]���� �3K�m��{� ?jGO(��l�6ˑQ������!eJ���I�jg!�W/yvz���c�K�~�pQ��fc�we�74ƽ���B��8�N��:��p���%+�Z��^ֆTw{<�����VW����l�C�L3�:��-3�8��s��.-:�� 3q
<E���;��;�7�x�?_���å'�~Jwy}��0�8RM��kJ�5�f��F�	0IH#7E�ߤ$ 8�-�C7�����.Z��jv�q1��3;IZp����=�j~�7%� ������fU�뗍'�@�zA�M�^k�-���[?�ePB���*�v̜T�*?L�q��r���|�p���H���#��pGZ�/r�ɘ�lL����r�,�1Ӿ���-֩����O���?��w�vsa�}��۵��7b��~����	X�H�������'�p��nQ�ÇR2#:��f���ꨆ��l��8X$m��E{��C@�>Wg
�j^�R�����_S��u�q�Xm�C)$JE�gP�V�:V߿=P�s���#:q�1l���X)H@�2)��x����ǳ����E�;����ߵU�4�fW����/E�R�]%����:K�t�c	��^t���l�«���xnR��6�^2���/�6&���U3��2#TjT6�L
5l��W�u�^h��B����eR?���m�:�%>��݇��PJFʦ��_��k�n�G��Cm۟��S��ޭ;�V$���4xR��(L4ĝ�b��=��.�}O�``A||���!��`�ܮ��X��&��QG��TsJ�a7��$_�5.L�\D��?_��lV��z���!{OW�R��y��U4s�b�=�֑W`�8v��4?,�y$k�jۀ��5f|����f�'��744n>PȬT��� �������Z�J䂠@�}���k�c{3������M��a���d�'��ӥ ��6�J�'������ۜ���r`������n)�����ٶ�a��R�/"�H_	xs��)�$��Q��+QlDs�þ�a=V{g��$)}�<F���({g�j�g{#�]�ͽ=�M^��|&C<�NO����1F�ch��R�����Q� �K-/�U�Y ����y�n���>6�s�A��$��Ot3-Şs/]Ж���4'�呈�sJ�s4[��'��\�Bw��h��j:���ܾCC/��h\V��:���A��²U:F������i_9��0��;�����U��^����ٛq,�6�si��u��,I�	�/�q��-N+q��L�h6��5���\��E��ͼ*=	�g��oP��_����!�4*��R2�$��gN���Q� ��P�uf[�:�&�Yc$ۀܿ�+�ăo��@����ei�*Z�Ƨ�����j�k�O)M�Ơy��P<F��e?ٗ%#�V�"��--�~L��u��ۘ���"����r?��.Fv��<@�!SI���f�}��k���sf��������E�[l�oqۢd��:��1bi�n	���)� H�ƺ�B���� ����G{>����*��R�q��5RH��[2���'�Y�ZB��
 �4�s6�_��	�_�Մ}S���3uH��#v��ewĨ��,�`)�Ƙ^5��8=�Tz�V؈�	�Mzf�y:�#�� �w̹���m����P�8�;����B�qW~8__��]��L�S��̐�wotv�%ͼ�i_�y�%,�J�����(���7H�rSW�RS����ՠ��Y��u��?�o�Zx4�4�y���5�1�6O�����F�����_+z�xM<R?����IS<R����3�����踲��� (���F����l9外<)#�unٕ C�{��N-|.=��l�( _��AA�r���AÍ�_o��>��b��OÇ�Ű(�u���*Z��ߠC;˰�s�Tq[M@�Ѳ���WǊ�Bk��w�[i��&��7��`?��r�a��]�y�<?���]�(�>2T)�+ٷQZw$D��VP���5B=�G�/KSa�/�����6��L���̚�˥��N�el��*�kyܕ��/�jFY �.��܎��÷4ZQ�Uu�G�l�@�t��@�l�@�s0zL��
�r�JZAOJ�j%��-��V��?K)-��'����絽Z���I!���P<A��l!��Ȯ*���U�T�?���	�`���s��k�nO��i�#����bI�D��\a׼l����
�+�&�W�*5���Ɵy5��Z�Tb�e���f�����LZx�ހ<5�5	���
��/�h߲�Vׂ�M�Z��U��
���ώ���ӊ9����aߡ��ݺW�;���)%-�u�n}�'�!V���V 8�:�B���� Y==�v!H�a�{��9�^(D��P�F0��8��I?�,�w�ƒ\��8Z�}U8ҡ�O��t����b��]	JF��}�􋿗K�P�ld7w	Q�W*y㠔��\��W�LF�a��\�u�!4�x�1/�@��/���{�u��,�)���wЪt8j��{0z����*	��m�&i �L�1�K��hS����������?�l�N��^���́�~�P5H��=a�刿�g�o/���#��L��� J��z`/>R�/l/�9|$P(�z%w��8*������#-O�Xp�a!��;W�!�W�0q����H;w���ӕ�G�u��k���ޒzT�S�Q�KA����8�DP#���8❦c�o<��Ly�]_�6ӿ<��_&�fH�_�ټN����2�d3�TK��ڌ]����vG��ә��C��-X��]8���|�n-�f^�x
�s߅������h�] 2��$���s>~����"Kԉ�kr�1�PQ	���:��U���3�7���|�X�@��2��k��t��8���5�j���%���f>S�=8����(q#������oz&b$����=i�\��!���(������H�Z={���+�M�\�R��{��Ơ��^�#M��#.��/Z��]&�=hl���2�U����=������سX�2n�m�a���?��ҎO�a�����+3_n��2��Dt�>B�`~�$�o�ͯ��}�d]��96ɧN��$�f|�������N��B��u��"�ɒ?��:@.�x�jِ�.�܏l��d.��W%B��<UwK%d�U\M���R
��GKZ��_4�ԕ���>��ivM!�y�4)d(|}�z_�����������o(�CJ�?�<TJ1�� T9��Y�r{&�Ǵ���˧^Wtc�m�!�<�.!��yY<���C��+�45��SV�ex�NmA1S�_�[{k)���[�,�zr�M���x��0�y�q� DV8�$���M��`_p	��3���U ��D��O#��FQ�:�q��n��7)S�e9zG�ɟ.� �1MMQx��^����8�=O$N�{(uW�?+��涗�`Y���6�3$;~���"t���\�^�)�쑰Il��2Rl����@v"����Kǥ�wb~>V��� ��� SP�
��jĀ��М9�ʨ�{1����+�n9��]�ޞ1�&Xb^�М��b)�-~���س�VmLgBK}��]m��7J����Ĥ��l>J�L@�'O��׳/�& ���z�D�?�A��d�v!Y{�࣒(�߈<鱲2v���_K,)�{ud���
�,aeĐ�n�������Uӎ\$�r%�E�	��Y��"D��M��$n������ˑș���1 �K4@�\1�(�З�7����.9BI	{3�J�4[�^��t�B�N��H_��}�M#y8�<�50EJ��%7�6ji���KC̓@�3�2�v�I���TX	V}�PT$Qg�]n������Ь��ъ}��g(��o,�SB�4�k������4Y�c�Y������ې��D�u&@��=��=;�>~�!��dS�D�xrT�0�[�rM�[�}���\�+O�����[���[*G:��`Le�:=���������Ӓ�=������< ��<�E�L^��.���0ω�k�����vB�V�|��S[P~�~.�VI��7cC�4>����]��nH��kJ��v�2�Z�zk� ��ȆZ�6`��W#Yl����{��j��1%�$�_�#Rh%k��fW��	��\w�(}1��h� 6�6ԭS��+�� ���.��zQ@��u<�Ϊ��R�5�����g���oڠ�`��a5.���	�F�W�������� �Y�n�<i�QR!�٢�sTx�|���E�ǿ�g��G��M��X(�����Q��~�AbRJ�a�SlN�{�J'%SS���5O�-�רɉZ�����7��ڟu6��q"$<K7�L�MebϟrA�����ǵ��~ة�H(��+���@�(II0�Ȅ��������Jf���9̾��k�'��N�w���39�p9;�l����ɨ�XWܼ�����&*�ٮ0�u@X�W�n���h����0��ؖ�\H����/I�+������]ܤx�>��1�Aչ?�|���Z����Y�p-� W ;`V�&�������{������]pFG@Ok3�Fj�'"g�`%B<41����V��?�b���a59��i�|�M�=�dc��D��s�m���h$W�]~IyPѺ����4�R�o}�1�ry;�r�7/x��p`��-���ޭxT���68����ߐ�
���j5@Ta9WZ��@�g�~\�5��ҽ�t���b�69l0/��ı.K[�#���vi��C��	o�~�6L���&M�Cq���n�q�"G\nȎ|�t�-k�@A��N�[=R�z.����}QV2��Q�(4ҋt-��������T&����NJ͹����f��iQ������#�7?�(�zh��Q�Q��p`}d%z�H>ñ��0��7�@Y�}�Wu]/fѕ�?����c@�	q\x�߀��'K�(�6�������7��E9�=�셸�.����S�;�%�X�j�p����4�ߑy�������B[`����끰�bng�+9P��~���*/oP4,3�b�&�Ԫ�%;��kT�.� .����n�6I���I�c$X�߬�-|�k���_� ���w�+������?�`�0�B�c�������&�������������vT=�:7a�]�c� �$�syQsZ�T�՗Hu+��F�+F�,x�BÅI*,�O�{���Z���:�w����~��Hd��%1��כ!��؇�՗?�>���=&U�P��oZ�2m!��ҷ�'�D���36���Flug�_�Ã�u�`�8#�4^0�=-���z"	����d�޵��x�#���:�Km렢������1w��t��9�G�O^*i��#���M���j�#'��K��*�G�hT'7?��#G�-x,����L�����V�_7��������q�TQ���=�"��aQ���GwV=Q�D�6�1��]�=M�a�'S�Ac���d�0�fK�~����$ml��ý��癙���$}�Y�*T�������kl+<K�L�C\7�F���e�Yg*s,��^���i[�X�; �Q������o���(ŷX�o�4ՎL��Q$�JM2P&n�bt���>;�Z��z��el�P�i�Xc�L�j�ۏ��EU��&@%��A�%F�zCܐq���A�����pK���e�wP�.�z/@5�8rd�� �M����0�$p�B�� �!����.,��@k�.<�Yz�fu7���<��m0�5w����h�A�t��0���=�� lu�z���s��lq	G���_Q��x�kc-G~i&<������1Y"���.��Iޟ0����	�aK�_��^��@j�\c��X� �ʿ|@R�qC�����}�'�ͦr�T-p�񽼓^ӌ���W�`4��@�q��%�:]���7���{�i�*T�d��u��I��_<�g����C�s�I4`؃9Ҙ�Oc����Ǣ fw���7k���l�M.)]��:h�2�oŤ���yR��q0|qV'\�K�U&Ƶ�� {���Sj����0�S��o�/�82Sn�8]*M��ؑ��u6�'�V����P2C�ڔI)t���dJs-����E�W���o2x�+�>��s��Qհ3Е{\�I*��e�b�t�Z-�r�؆Ʊu���&�'�3Cͯ �U�@�#��m����;�>��� ��:���6�u����������aa���;!n �"�l�Y5�T���/\i �  {_H����mĀ_�D_w�q�[�`{Fw�\�ޱ?X(#��J�h��ڷ��ct�S�K�]v��@,D�>,"���A_Ʀ�J�~z����3b�S�L��8�g۵�I��^���0R�C42�C�����eF�Y0b��L��W��j	&�!��B�cZ	z;Cl?�|Fm;�ڱ���
�� F�	L�[_�}Zc"$���=������v��f�i�FJ�q��M�Ñ5g��7xAx\UV��Q-b�� w�C@*��l鄍ד!�;Ah���Vʸ�T�����	���r���^�~�f2�)s���C>V�)\XKfy��EI�Ђ�Ot�������!���i��$N0.��������g��;���JH�����>lM>� ��D� ��J��ۆ�fNa�V�5[+�w��W�iV��3G�����J���4E�||����9O�C��T�׏���-2A��l=�ͪ!������t$]��a��4�xK�L��)[�#��4��3!R�|i��8��Ɨ֍Mآ` r@�X��󷬤��i�a:�&
<������s�'�d��P���k+Կ  ��qtTz��)i�߁3	���1��L�C]��E����� ���6fm�k���s�a?���'�_��ӜweE��'��+���bOo!Fн�ꬍT��8[9T��Eʷ��2�I$���V'�DU}+d�~q��.$�'��LKsU�%�;�$q�@�;�:{"XWIk��r��_��8�cc���ճkV#L���N��{�I��f\����ʠ����[���>+s����d5�c�O��l�7M���>���uc�Qe~�R��n���܃�8������#5�[���j'�ڍ��;��\wsV �C�-�
I��.x�){e�0�\˨�Yx3��x1R�+��*�h�1C�O�ma�	�Ww�`�}���r�s����5w&�_Cx�n$�1"�`�+CӇtŏ�n��<:d8�U�*d.�I���U��k+<%����e�hR��CCjtZ�|�uUZ���G�3�8��/y<F�=*;�=U��LsTz���w�h%�T�����U�P�q�c�.Ҵ1��L8��9�����,��;�6�^h�0��0�jsl�V �N�5Ϧ���*g(~U��7V	�cD��O�N	5�VÑ�g�t(�>r�D9 �G|�ŝ"��r\�ށD�Z�)*	�� R�Xĭ�*����wm&�V���W=���3��X�����
���v���\�@�V���7v�K��	X���z}|�@�B�tm�����T�m<A��&;�~��'G��7����]�9N��@�V�kZ#�JV��;+"����q����f+.{���l�\�����E��^��m͆`��Z�1����bx5���Sw\f�s�/����z������ۋ�bR���alrO#�l�y�iVwߠ
Q̓�7�@��B��HM-��Y�%\k��Zצt�J��%��= :��̲��F�a��?'򑝯������޾6�֌�����^ƾ��X`vV�!�hM:��-}�3:���U�xpO"�}���f�v�.�0��W��U5)K��M"�Q�Zm"
}tz�u��ߤ�&|	����k��3FQ�ޫ�����:Q5���(y�*ɲ��j��s���e$���[*���j�\ax��V@�=�b�˗]j����l�����a�QSq\�@St�����2I���.k=������?���>EC¨���RY4a�j@Z9��>B�Pv����փ-��Kέcu�HfѺ:q�:ݼ�;[�ᖙ�Ӹ|�f���U�.��Vn0[8��*���H�9B���`nod��IF'��ݷ��֎���P�Tg�C5��\S;�������v��M����X���.�d���=L��I��|�Q�Z�>���Nj�E��#A[�PS���?Ŧ����Ѽ�˽qy5�����*��F��!,�U�͙��6"��� �pnk�~��,�Cߚ�\��J�\H�@���z*�!X���MyR�ai�����]�M���U����L�M�D3tL&
)0���I����E�x	�''۾�d�o�0�� ��I��SQ�����N�5�k�ZN�!�$\��\a�S�vl��k	*#�:���i9"!�>��X��(��.q��_��t��_Q>�ʗÛJ+�LtN��V���8tӋ��*�bs4fR�h.�#U�̄5��_�qA��I+Vy����43.Z��不q��v��f�,hA`��֒S�64�6���� �څX,�~?u��^����h��(Sk�X#��S?�7<��2��H�!���� �����Hf�#�&�%�Jq��؀����`���*1\_�r�2�)�M\��5I�1�]���C-��5�\fY.��.��2Ť��^�������-B\`Aƣ���ȖG�	2����4�G�C����{��#��&y	����plq�3���#�kP�Ӡ�
Q`�f��y`�kKz�L@6�V��������y545T&����i��d	������ڼ�s�n���U�b!�+έv���~��6�6���wԚ��!�l>������z�~�_щ;�!��m��J�s�]�����PX7�|:�����^��_Q�;��]��h��<����S ��xt����~Zy!o��??ÖL��4�k	�.J���(��#�K�����-��$�EB(o�m��\OT�L�ck��$���	D��Zu�ɭu׮{���@h�ceƟ���C�hU���
6��h詭_�W��~WD�r���b�x�.��x'&.�P<!���Fi"Ake��h1G�&���r�9"��/�ݜӲHJl��cJ R�&�ĕ��E8k����^���6En��޼Ayj&��y�@:Do%�(-}$�*]�oc��9jvg��-5�%�g�
��肊4�]Z)�$ӹkBXO��o�з�ŒnL�n��=�c��bEq������PЃ�-p����wȧ���?��6�I��_��y�u����"؄W6j�a���	BWS5����#�f�0��wf�Qsp݄�C�`N�:���-6�C@�v܇Ke�	���!��n�}��.!�)����;���@�9�:�6�<�|�Toö9�|*�}wW�-k����_��=-�h��˽����G=�1p"�s���j�3��v�N�N�U(^�Zz~{������֬AO����R��C�q ��Ss��9��c�狁��e�	U�s� ��Y�Z���I3��!g�?�;kLDZF��k�ZZ�N;yP,�ާ𠷧��p��E�*���Nm�×$��5��V��	�v��ڌN���c-8���؆yr����%�Q2i�7e�oM��֎�ZA=wz%c�����:�IPoN4���)5���E��T��s���-��)(7�j�!�����s*/O԰�rm�y4E�8 ��������L�NDI���vWD)�!Jq�D[�9W���?���`���P���If-e��k汯�G�GG�y�w.x���uj��O�a�������G�Lp��`���	j9c�=zi(g���d���4/�O���_δ����<�5#)�0�V�|/#�  $Z����p�[���S�4ЀB�hu�聋�����`䦿�6��p����#g�ȿ�@�)1�N7�SO�̻���%;^*_�?������{s���9��k�\���us8bV4߀�<J8ET���0E9/I��3�O뫓b�)XO��G��`:��v�"a�0EAf�L�Gj¸)�͊�#w�i���P��".P�ظچ����	�|��G������k�d�7˭>V!䓏�諐u��g-������@��J)����eVR�}I]�s8��+6邑(mtKם�c�)bc��Pd#H��k%�
m�1���Ť�`�Y�"��g��V�����f?�v�W=)0f4D'û8��t�e����֧�E�uF�����suJk:�������E��_j6ǳ9
�ȕ��Ѝ��Ae �^>fH;��A�Zl�M���[Ȗ纪�xӆ8Y�ے<�S�\v4*g����RѤ�k1ӝ]I4F�H	f˚m�7Ad�8'�1 P�z�`�:���J�3*e��&U����΂0dIt�X�3,LNi�z�wUjp��O!%���%F�����;��}���\��A	�ˈ�l�*���[Qrv�V�bJ���J� �	�j!��Y�Xe:�;:,o�/�x��Q3��ͣ��٩l$W7���,H,1~eo3��M`�.[�,�!���}�?
�>@��O{�����`��o�������ܔc��1��O�P��(ϛ���w����ZoKҚO�+�B��ᆧR��7�����p'�#�we�}��xi�4�ר�Nʸe�N��u{�[��tr�~�񶉔�Ni�����ټ0	^�x:���k�w#(�P��_�Tl��>	�h 1��	8G=�XT@ڶ=	I��mB�l����Hl�O"@�q?H���2-�R"� ��H�5S�`�m�-k���Y7�N�GX!^@��y
�}�J�G���7t���t��S��֑?��r,�Rp1�:C}e4B˪C��d�W��i�Z��<d`CYBohӊp?�
 l&T��~�&�seT�K�l�Uͣt�]��;F&�jv��aՀRȊ/6zp�&W��y��7�bQ��݇0��^��9�,�-p�n'���ǽx!6+������w�y�����;��LAO���}�;�ix�c��o^���k�޽�2tM�8�.7�x����&���҈ j�=ns�#�I����5ZV0�r�Gz�����5I�t�N_�J��x�b_�d��S3�a�f>oS�1�)�;h��%����x���v�����P��L5�����3����ہO�8�U��Tt�l)��F�0�9K'����U=��
�[4��8G�Ό`�ݕ�t��Z�(��UG���Rt8�9�*���=<��(�6Sҥ�b��+/oYU�'-� ��(X�:�� �m�b�A"9}���E������Ru3y>(�щs�4}֏�p��e��?�%g�꣬Ϩ�35���cz= G�5G��ɷ��zsT��Z]�ZltG���n�t.�a���1E�=��t��d��OvI�'�x�#+HY\���"��S������nK����;�A����J��-��m!��(�_��āWP�#��VwS9R��t�^��4W ���tl�z�g���k�U^&O�(�l�x�������<�B�z���t[�pX۴�$�6i1=o1����G�����/g#���lMXp�'v�.����	����S���`�԰�j߁{�NU��ࠜp'�3��.�|�xr)�$1b?��Ͱ� V3�5�Y8X�!e�>v�_3rZ���C�G�֥�`��mi^l)6Z��`��xtf�G>n7�n�m�������K�S*����Ba�xqʁ���'k@�I������]�ڼj��MI���]<u�5��J�Տ@ ����c���1#�S���\��V*�5�@��
M��J �$@����u� ��=����,��ւ��}bׅ�t��C×���}�s��b
 pS12%q�1��Y_{8�3��c��l�H��&]��>�|97D� #��rA���Q�e���v�kH���l�Ѥ#ǸX-Cs,�oؖ���z`�$��<�zi��oV[j���S��)ְ��Q~����㜀���I��PA���إ1f��;�~�@PJ�Z�� �3�t�88�=���ǘ��r�ċu��`�n�k��G��(�h���Uv�����J��/��.�o+�lO��2]��A]�x5:�����6
���Te��AF�?��*�07a����,�^��5X�kS���KA:��<e�r��( ��Q��>��B��E�ܦ�iwX��M�l�W���RR*�#�J(ɻv4�����<�����J�g|���E���Q�*����Qu�$�^�R�O�e�_b���W�}��V�W`�T=�c�o�+�M<�6.d��GrGwc�u��*v�֦�{/�y���\��Iѻ?븪-�٩~`��.��z��A�bu*��kQTt˜@C /�e�*0��f��GlY�%+�{��M.��n�#���RW=zHX��$�@<��g��&OZA��]�3Xܐ�#���IśG����$4V�)���W�qa���!��W؝�-��(i	�#��$��?wGT�ԧ��}���^@>�V��������2�L�I����W�/"��@���TQ�Ą�� '�ЏK�3����q�N\��m�J��&��G�Z@{S�m����#�� :w�&J�0+�;�;�Xa�;�7%$�@��Z��1b��U�Z@��'y���&Tf���Lv��Ld'�W��>���*0�?r�=�z; ��|��l'LI��K���u����U_v!6��\�ܥ+l׿��B�V�	?*�r��b�*����p�)Pi2`��fd����%*�b�!���9���E�{$��ĜV���(H[�o"f�A��N]J`Eޑ�D�O�'�ޓh��(va2��]��T�|M��9Y�p;f��	�X]u�zg�h>_�աpdq{�"rd�������T:ĚZ�|��L-d'x�f���Ϳ���$ �4% 5�kG��3�L� ���x��]ϼW�!"����=��х&����~ö�V5AM�xX8]*���ۻ@�Fb�%ae|��ސ����1��ＵV�@���<m��B��>��}H��A� G��*���vr�-�Qk�_<���t��6܋2\4���M����9�i�4�=�R�����-/�(>����C�R�ߨ<�����N�ӄ 7����Z��1ίݟ��7��2I���Q�XrF{�6@�p,���Q��e:{V��	Eʪ;�:w��ɰo��E%���|y����k���+��C��G�@&}���MR�M=��ni�N�쬂�:ː���d|���֢j���5b��������
Wo����<#X�i�c&���L2ʯ��2op.��1d�ٰ"��±�F���Wb
��``�WC��E��\��o��2�Ş�`��-G��"�T#9�T���ra]E�Ɂ�}8(Q{vK�y������|?���)雳��)2�8�貍돌�7zi�I��b]���8H7j�]�-�[ݙ�'��,̀q�tNh�Wʩ��n6�aIJT:f��V;�Y��m�a�e}n��Hj���nK ��� ל���!�0����._4gt),�z(�6���p>E����xhL	�RE�+֍�2A�	��p�HZb�/��xE���aB�a�c9�r9(h��I�IKN6����q_��JLI{��؆V�d#LA+�ߟ�@yub""t����F���B���v��K�)�4��r9R0'��X+\n9[�b���cPa�k�A�E�t8����5�;����v^W�z~V�iN������z͒��+��C@��P����t�ƻ�	�|z�AE?��ʶ�>����2V��O��2�� �7C�l&O%b�n�0¢&��M�w�o<��v �0ȥm@}�$��n(h���p�c�F�n޵E"i*e�O��[�S���\�F�wp��1�H/�_���r'�-/���Jw�:x_��s�ꈿkgZ�i���ECC���%��m��k�y@��4�O�AJt��v�*#�Y25�#��ɮ���ʥ5���_�/A�yR#5^�[�#9���i�� ��AƓaN}g��^�i��ku�P�V�~�GwJ�~�ϓ��uЯ�\a�sU��9Ԧte��BB]C�w1U��y2�Z-w����3b�.��`�΂ �ӹ=Ţ@P�	 m����MRϾ[{q���Č31��!s	`�Dn9��ٗ�hdlZ�����utw���w+���6{f�O�u�ܨu�8(c`�w4�w.T�Lgh�2�Ri;��wX�Q����ck�bCh�"�Y�6���S��z�ԗ=uK~�X�}/������RG�_���}s?�T�F6E�W�X �Ң�K�G������.�e!�l��Go���Y��r�\_0<2{�q��
��{X�!�ݰz����rEg�wiݷ���5���ff���X�h>}�9a�B�)�d$/<�[��pf5�vw�B��S�	�k��*���?R
.D�d��b;��h_o�����-��R8�tsi����h�k0i����G���[��hC�D8���i�UO���-�yXo�����W�pT;�8��P�_���n�O��!�V�����<2�6n�^�^��XЬ�{��~C8k��ics�D�����؞�	^� �H��bꙀ0,5�Fɷ�Q�!ԕ����$�G�c6���ݍq/Ŭ���`�@�{�~�?�����j��o��p��@��}����NЪK1�Li��s�̚��k�z��=�\vC����H�V�(��~�JDa���D[�WEb+o��o���q��C)-���t��C�q��:[�[�H�S.W0��,_�
-X���P:D�HE�w�R�ƛC�<˼t�S��Djyx�!N�d
��ܥ�J��L�+<)!kp8{�2��H��x�֋_X�'oRTk��t�N����Q�M}���%���-��7�MGY�-f\�����g�OҀ�Xp@�柜��g~������_�T�=�{#�I$�j��W���q����{߉plT��$ɫ��K���{H���Q����őX��T�Ձ%K�QM��wΡ�`K�i���h?���s���7�TE���
c/=��G,W��!D��KCH9ƭ�u���f�ރlW��mw-e�+N����#��{�69g6��_A9�_[����"�;������I���5q�1�QD���"�{�AY���"/ =Tc��<>*�WWR��N�hz%h���T����?��TJ�K�*����1Sy[���k^�Y'���`B��(Gt!|��X�)m�9��x��A������;$'-Q>r�ɱ�/~�h�.R�'�^��zmx׶�1a���c��� 	yjjF����ˋ��[��i�F����4�����:) �V݋V�0���"3� y!S8h�y�*�f��0"m��iZt'��qrZ��;�B]����cJ�<@v-��سpsF��3Rk��	�0ؿ��lF�a��M:��0���	P妲�=�t1����B|�����^�H���؁���m�}�K@�ް�8�D���`���(�FV��r I����u��Z��MF��puz�����G#�#(��-�*��|�Z�lDf*�H"*��{�����C�xա(��o��\���>�8�VCye
mt!B��k��o]��ٌey�U�ؙv)x3{�[��K���!�8��}*%&Ry�u��I������n�NR)u�_;U����G�qk�~��Q뢻d@�ɂ��������À;�B��f%gߤ��ZC��)qՅ���ssg(���'E�R�R��a�F)'/�OcK'3]��g0)NBhk@����{�e�������
������ �������0j��_L��E�����~��	n8��jP��p�(N��àkOM\8��qn )@�W�����'G�?Ťw2:TF�O�<;uW�H��<��:�D��Awogl����yj W��椡�}��"G���x%�?�6�GiF�n� �Y�kr���I_}�{i��<(���Gna�b6�*���?WQdB���I��I;�ީԟ�2����L1]?�⮷)��E��s��� �W`��U%�G�=Gs�Y�9:An2S��P�o���0v�6� �u,���Q�}�9$� �JB�Ȭ��K/t	��B"mH��%��P���oN$��;�ްQ��z�X��)�1G���ڲ�:3�ki����p(vtMAN�L�ԁZ)�4�N�W�S;ŕ�>ޕ�b�Ҫx�����t f�y}�S��F�N����Y��{�*��ˬv�M&r�U�/��3�L�\2-Sll�� X+z�ԙ7Ĩ�@�F}��7낦�ߟ��fQR����je��ｅ�r?��Ob����w�O�,�ϣ���2�d㔓a���P�&�e>�$���t���`���&<������K�诨R�С8��	@�����i�F�@ �R�����ʯ�Ch��~rqfs�q���m�lD�R1&�S䫊g-���]?bi1��$	��:�_f�du��Ȫr���&D@���ё�� VE�pY��~g1�ݝ�������ϥ�}A���u���M(!�ťd��#;vN�u��&`C*���ъ��ɲ���U)ވn�6C���qgo�Y��C���B���]؎��x�;�ھ�kV�PI��u�����o�6��f�����鹻�����䟦$;fww�e�d�)K�Q3��$P��b�����hr+�9^�"�U�3-$W����[���G�q��9�H��њG`ُ|�[���0�;�$��Wp�u\;Ȥ��bl�9��z��*��m������]�f���i���m�3�@���_����3n~78� |���ב�}�P�^���-�d��lZ���1nS�����wW�s�ǐ�;��W�6��;U�$�s����_�:`�U?�-p�f\½ù��ͅ�E���M4{R����s�eP�Ihh'7��9��W�K���\7�g�JA�f�N{��S6v�� ;U��0\��Y��7���O.��C �,]�i�:(��ch3j%�`0T�Ҍ�O�y X�%����/r���'�3ST:)��2�(���^�bͬ�1K�D�{�K\�ub����\�&c痲�Ł.Q[��	:��կ)�͎Db���y;�fhQ�����T�Z y#��ۆ<%�}��D���di���đ�Q���^�k�$n�Ptab�W��+Ċ��O>4�E��j�:�{�[3���W�F�*����l�Ԧ��(e�Y�I����7ս���qL�ہF��@�5#��+[N	�~C��J���8����f������HhRC����?z�%��7v<X��t�*�J�זK��妾�L �����H�qn�L�Q�7,��A��jXm~��>5�b����	�An�ֈ�J(�'uN�r�X��"=4&���]v��'�r=���*���n�7�}1~��خ�b���;��F�� ����Y5e�Pc(���(�e�< x��fgZ|��2!4>��.�;�d����.�]�
�&��7���3Q3J��a�Lm��ʤ����|e>c|[�r?mv�߅i��Z�w�<�<۟ήf[=F��J�D4�����e��_�,7Ntu��!��՜Ȝ�N�l�HEh����jS�z�ើ�^�9��d[�
L�s�U��Fe �d�QB�@;7_>OZq�=������c�=�M��.]�Ȥց�@w�"�G\>��^l���7��R�صF�F��֫���<�i�����:BG2�W�bC��:�q_��;�QȠ*a�����=�<�<���,�X�p��9�����G%�����R�z-�"�雪[��'�1<���-D�ڭ�>��L���g1̚��t�lAt���,Rce�^��>�����h�͉�ű���G:9ͱ�������z�S/e�\R4��W�Fw��	@\�V ����cv�༧�d�����]�d;�ƿM��G�QiqLR�N�e}
�ƶsϨ�D&�(&.��&�jM�gP��=2���w������<��q�*��	y�*��Z҂, ����a��z֨���@�F;�ѻQ޸�u7��*l	�t"b�gfK6��{����9�1m�ikv�w�%��
����Hj���Jұ����T8j�8�h���{�x%���l} �^̐��&�F��ʴ����eW��F��t����;�]T��T�.���-��>̅�9�/����{y���W�JH5xAD�+Ai֏��+���R�}5����bl�{��m3�f:���C��	,��=O/�7�3�(��W���t��ܡA�i����1�JR��J�R��؋Q��ug��*XU/	��_�naz�r1�1ߪ	h�`�P�FQbǛ*A�`�5#r4vm�[S�a��`Ɓ�L�8����$���$W�M�"���1�l��u§�"p�&����l��-�B��+��@��b�9�݉IGB�u��i����~dqQ>�dC3
�'����?A��şx@D�mԹ8k��a�첥f��.���/�F���`�'���WIGJ: �b`��|)�
r���5c��NOtp��o�0��X��	h��v`8q[fR�5e^�R�Y�rO����`"�a0Qa��ǀ��гr���ǗX�V����:�C���捭���X$��sZ����{��V}��Χ�_))+�}1d�?L�?4����z��.��j����UF/�[�AXG����\�;�x/yh�>f�N;{0�����H���8�fj�9w0p�h�+_������	�o�U�����[IM(��M��g��t!���aY3��cf2�&��/��΄ώA���\`����}f�d��M-$�"�RO0&��ly`��s��E]W7DSevN�OW]y���E�n�h�O��{yHy�P6͡hQ="�������$8u7����?ܭ��	-Y����r���y���{�?�++�v��Gj�+,�$�L�q��y�Lb�7𣤁���,{��\���_q(���\����
=��f+�7��	�=�X�6+����p��'枖9�pC�j���l%$����T�h�єQ��v\q�y����^�D ~ps���Ue���*�p��AѰ0;��$L�{�6������}e�hߏ���-M�^���F��2E�H���_��<�:�C>�{Κ�RUW��"V�Z>\��|�e��8�'��1�i河sx���̅D��31�-�8|Ҽ^���iZ��(��O��$̗��R/4��a�OX�J
�XIe���Zpu|M-�IMKҦw��O�9�`p�d�������r�@M	[�%*�������:�&	ح�5o�F������D��"���F �\LQb-���+��N�3�C��n����"2�.�Α��"^ ����5<9|Ui�L�$ٔ�w��Q9�bc5/f֨n������ߟ����[��~}:5]��ku�]���ky#�<jH=F���`=(�L�]2/s�KՕ������7����`%�`�G:��͚/���(8��A^��?��l�SW(�o�Wpe^�B$�0�k`Ek�����&�u:2Ƅ����k��uTMc��m��:�����H��X/Tم7�Z����尨�  P�6�}Sa!��똣���c�ժ�4'	�b�́���6D�����B��G�N����=��Rg��ӊ�Я�
���f�����EE̶)��m*��%������/�Ҽ<M�����i�8 ~���D���x�&�Sl�� aT?���X'��k��)E�������ٝBMXD�>�}S<�Ƈ_���֤W��zeZ{<Ŏ�㲹w�����)0��f9����|s,_ȿ(o�����xq8Y�/�m�E �(�m_J'0,ܱ�҈�A���mS[���}ڇ�B�{�92�B�4>L�hӬ'�[���X�T��=�fldS���q�#��J�����#ǖF�#���@CU�iJ��x7ͳp�>D��Z�O[��*�)�Hb�@i���d�T.�����!:+��x�j ����?�fܔ��l��%'..���PJ���jޘ)��d�k��Rm��ib�ڱ�V@��Q�.��ki���~< ?;�
j���_�Г����f�_C�«�'(��-��Ĉ��+U{��@,=�6B�t�dBX�'�}r�c_��آ�Yʷ�,@�l�	^@��`gQt9rk����2ܧ�S�Ơ[�#�Gf��iZ�'���n��a�������A?��-��z�)f�x??$a�������>?"�]e�A�Q��d�K.�I��ZWZ1��+#��I��ϩ��_��N�,j��=�lS��ECgBJ�B7�%�7��xX[U3�ْ��i�pA�!�Y�Ͻnl�8c�M=���qk��H_�;SH�@��=�Ug5F,M��ׁ(���	 x�ߍ���O ���rK������ז���,��&|�u6�%�W�����h���o�>�2�;Rs[�6V��]=��{adS󃓰hU�6���G4�
ϡ��实��1Jp��6X����'{}w��g�gG� �x�Z&��0�@�����lE1m��������?Rw��q�꧘#��m��
�Ӻ���٩r�vj%���Z>���zW�g~PӅl���P��|��������00��Cf��}K,΢�����Q�!hm#2 ����~���d�+�dL�>�i���n�#�k:1���*`)RzG�q$��/��`B"i�A;�:��ՠY�<�-��Ǎ�Xq��A8��A��Gy��B*\V��3;���i����o�G1��Q����%�<:u�%U���\�Z���3���� ��p�pI������m��!�Yr�W��Õ
D��ɁQ�х��G�`?C�%���"�D[�!��I�9zpL�9#dKQ�����_j~"���#�KJ]~���I��E�/�:j�:[���bō2lm�ֿ��8z���yz��ހ���<^u��d>$9�F�	�A��l]R�I�h�e�B�z^F,�!6ƝS�tK=�����^�j5a�8y��c�x]��	�V���2uka��F�1�qD7����������v� FYH�����U3JU�NN�jF38�iMg{h-<��jJ���u��1��'�I9�:�k��Qh��g��z�˭��v�v�D�9���RzXc|e�ż����#�R����)�<pP�k�x8Ǻ��I�ze�	��?���VK�!YZ��{V��D.��e����C�~��3����vo�G$����X?J�a����L<�\�>E����˚}���3%�c�]vz�����k���{h`�D�)v�e i���e3���و�VFv@����״�
��׎�����'�a�g̪��5�8.�'K��\+vb�|}�:GX�h<A�At�%I��K��|���f\q�İ����Hv�����EOJ�ǣ&��lS��[� -؀M�\T�ڋ
j��xT���}Ȗ�C�VwQ����K�맄�Nf�j�|r�{q�\DO��05�{h"p�W�NB3�xg�2��x���.���R�yjEB���@=V��U�e�? ��Ϙ�RZ���շ)�@mlq���Ļ�t�xV�c�_�����0Ȕ�B��˼0�cK��aw,�U�U9�L������Yt�g��'~NJ�dT������ۜ���aa�H�%�h��*�(3�C�Ķ���_>��^���}i�������ތ���~������\/�/���N�<{�a�N�2�x�5�8���o���������<��{���2c�,���u~S
�8��q�-���ТN�cVg���L�CJ6��-��R��\eăM̑־����~s!ORs&��p��km���1��1��K�pv+�v�����&�
#�ɱ�?#�P�w�e�mlʹߝ�F�`RI�%|-�m{�ѫ���U�#�t��% |�ݑd�B��6';�r��I_yR��E������ӵ�ҞP	�Vd����y#75��a1k�q��H���/��3���������?���ؔ�m���3�'��=",	�޽:���nt��奂�4tC��T1	���q"�¤\(a�	����!d��UK��(q'd�}H��� s�s������6��u'⻃h_5Hv����Bvp�K	4��t���L�cl�������5�j:".ՃY�7����s���ͪv�)��R$"˕*�A�'����`!��8}v�(��%�dr}V��Pȹ=����)�5�Ԓ;��Gvඍ۟""�P��&��1}�	b�p�4�8� ����Ru!��"�Տ"���)���&���$!TCi���	\�����1��t��V��f����i���iھ��6��&��u a�9~m�6"�lk�����=���BJ�߼S��l����{1�5d����C�=-+�r�����T�vQ2�N0Oצ���O0���1j$�������AFmUd��9ɉ���vE���a�e�y�~�t���$�`зd�k���zy�y©��8�V����J<xг�µ��н*�v�3�i���U 	��kxd��?1�� �IL]�bE�H�3"�qs� )~ �Ҁ<�ZJ�ed����ע"�W?�n�h^��+��h��k�A���02!\@��`�⢒:���-�Q�(�����z�3Q��q@�	 �`6��?	�C7{;�JN(ឫ��PGlj�Y������I�Gl=,�c
���	�A2����M%� lyLHrT YJR�]^�}�
$;�q���'�����'���}�f�̧_pt�-c_CMSﶯ���	R�9�*ςխyhT�n�Kez2�N��ܡ��r[��99~֕��h�L�+���9�IED����RUf?a�t�}�����⪾�p'87f���]���q�x^�c���Yy�����{ �Y���+�e�U�A[]�Z�;���j��;ٶ�U��#�:���idٵ�E U�[�����|4������%h��N2C��j�޶Q	P�Q3wwo��aJf�����>�1V�����`}V�����}>�I�0X��D����/"�Q&�wF�l���|o��,�jdO�i�8�H��[��4��j����9�\^�a���lh\?��2)��#��3�w�/����CC�y�}����&k�����qR�򙃯�B�f;�K�Տw�(�1����]�~���a�S<�y@e*�����R�YY@���8�	�eܑQ��&�`J-c���uE%�|o����Ժ�6��qW�}h!�����L����=���W��/�H�"�/�uwk���w4.w�5V�����D�5�r{��FIf�z1ύQ����G��HX�^�<�bR��@��DuU0�>鴎:���9f�RX��,�x�Z�Tz{(`� � s���z[Y��#�����$t�)}Լ��F�9޹fm1��pY/;�ܰ�l��JZ���\�k���U�o�dc�B�C9�O�����n?�|O��T*�Z����SCG_?����k�?�B����Vk'+��F�C�Ĵc:n�.VH����g2�J��h��t��7B�
�]4Us=D����k$��[�F�>ixa�q;��+[�}������Ֆs��&���թ)@�C`sh"��7;���;�'W�\����c7p����d�_	a�@%\��������l�BEؗr��>��.p��F�%)u���(�8d��⛃p&�m,��£s���)���*��`�,'���#+�Nv�ƜH���J�����D.��	sH}���ų��1���Ǘ��Q����+��(?��0/�.���T��3�EHFI��0HNjI��]����6�pM65~Q��k������l������]����䀴�뇥pa{����uZ�,#�nF�|0�����~��0�dD�q�i��F�ѱ�{�?Y��?�kQ�eh�ȸ6H!����|�e��(�:0����>I4:����^�d>�3�AaL����X3�� 0���?�,K�c:>G��Aө���
|�i��ڔ�r��v;��L?'ߡ�vd�e0{Y�f��_�LT��sV4�lv��Y�U�k���<@��q�>s+�R:�]�i�67K
k��K�5�������k���
�s*Š0V,7�Y�����x����0�����g���1����(ʐ���G�(ت*�Y��!����큺��A9DGp���qӠ�r�Wb[=����9q$��kz��#��D��+�t�ug�Y�8��T#���:P[y���������CY�iB��cbė��h�.�b�u�+Qks�4X�!e�VE|���`7q�|���#=trNDA����-��[|����ɨ��v)�\�\��4�tU;C&���r_Y29�Y���>�t�����z��PA�T���6A���E�����8%���uM-��q���@������O�cF�R�/��~����>r���k��K�h|Z�9��i���m�6:��J�z8ɮ���5�%ƌ�]>8��Q*�@/]�>�W^��*f�\�T�<�@���ME�Y*ޝԝ�a끚TΘN��3�IS1�2PyƤR��6(��g�o'(Z���P�J�������J%4jKo�g=Ʌ�}e��m>/+��:ш�HBh/�K�ا݇([X���'PXo-�o��ݕ�$h�����ǷW0�}X&kG��Jo���̈́?	F�C����?��e�"��
�����5$'ܯ@au�;����0p�Q���0��_��܅��+��w� [o:���/���e��c`Q��!�porP"�Pz-�������-�~�B�ff3-���!�������Zت7���Lg�܅Q{� ڪ7;��-�DV=Hd<�zC��K����b�Ũ��}�H!'3��$Jh@��z5����Cq��~f�V ����\��j�hx�.f`2b$�O��ĉ��\���=�'��Hm��ΫT�pZ��qq�<�I��#Vo���6���wJ�d�z�(�߉G#��v��ٔr��ydWǐ<�K��V�Bl���V����*��6斥\�XzC挳�i�2}N�/\'�RpZ��Y:�xƺ�lxoH�߂G��h8�ؗ��>3({� �Qꊛװ�𣷆�������A���v�_�e��Kp03�!߾��C�3\���F�0B=�����2��V��*�9���lh�/�$�\�U�懙a�ԗ�,;P���hKMX�ݕ���jW��q�B�zl��J�Q#�jnl}�,�f\�mw)(�l��ev<��G�
�u��.WCu�H�*�~� ���3�!�I}�Q��y�ڲE�/wV"��.x�Gj4ɿ#?K�"1�&0w�k����S�xl��B��VV0���v�qB�����0P���ɼ�j_�z��C�z���؏ܣ�dT�� ��Z���Ș��=�=��
*�g��4wu�^��o�U��-mI�.[)�~���H:�p�v	�UX��l.���9MBmH'��4�X����ƚ�_�[a��ae�I4�R�P�C��u��yS�YPI:�MƆd�B8����s�X^�w_�����#�:�fDA�R!�¢뺿� "Dq�cV��ٶ�$K���J`�����7��6�$���c���!���wswz<&="UQ��ח���;Єe=�͎0�*�Gm�E`�ÜF
����W���]�������xf-�6E�:&���FV�D�4�ŧ�T�;�e���¤݆�Q�Ƒz��`	q�W��@w���8��b�_��$�zd�)2� �=mi
������J��oK��F��[�o���F��-��֌�������q1ip�{�T��Q_՟��\~�yaU���۾ax0��N�{�#�uB�U����ߞhNU���GZ�3өwa�"|Da�g�ݞ�AE�W@��@{g�,Lg6ON%#��;I4��b{�����?ð��}�>݆�7sL��y���|c�����_M���E7���QuX
����8������]$]���4u�B��������C�R_3������]#�h���XX�����/WY�m���B|P:F���8�\?�V�y���@ ��JyI� $^�����K�t��|M�yw����S2�C+�����b&0�,�����Q��k��ĉ�$�����@ ��jniɑ�052v�����B�9���=����ű����?��L��vm���OBMz�w�K��q8mH�s�n�b!s�*��*����*�
h��j.BS��(6:q��VW��v>2��@�̞��AV���Q��4���z1�[�N�8p%������B��y���/(�zl��Esɏ[��:��E�2G=X�KS�6^�$.����������z�*"����ŏrz
������e��"yr�����h8�y�`�ly<>2sz��|����GB:P������l�QS�D�[�`^���_f] �<��fAʴ��I䃱4D����X���	��5����@���$����T�ffҎ�b�FҤ:Tc!j�v���fW�@��v�NM>�J�B��|.s�b"�}��`!��(?{�������j͒��b2]s�6>v�yƺ�&��-��)�Ay��@:�?G|����q�R�:�iDX`����� <���(��~.�Жz�S����sX/k�f����V�����!+����E7�S>�Q�%�����j�q�X|��+��Rh��< C�Ћ�����#.���t�r�e�Ā����?u���ѥ�m�2��[C���~ʄ��Uv^ ��҆ۈ�� �E
�R"���׺�%��ml�}�	-nFCo�:Ξ��N��5�ϔog��I�A��[$넢��k`v�SV����.H�����8������K�S��`X7r���v�G�0��|�|��8�V��-��/4xiֲsn
�����B�J��%��� \f��fs����Q<�⏗.���]:H�?���%l�L�:r�1^����I���Vg
�j�[+=�E��8��fV����P���o����#]A�;/Y�x0���W//�kI����Z���_���n�"�*��UZ��򉱄�wh|O��>���i����$�9EB�,R#�Nx���Q��������OR�CD��hKb_� ��.��X�I�,'��Þ�{`���m��JyT��k��I%�a�~��7n\˾��T�����5/pTT�1���\0/d1i�
䫘
��|Rn�/����2(�6,n��,ꪭy3�6NZ%��*h}��&���F�^2��bZ�~d���rF�D�?�r�-a����8��D��d�N\/@f��= ^/��}�X&9YV������/�.c��!�Y�U�����o-&O�z����#B��e�+Ѽ���~	\���+�����0�_���FveB�Lum;7yf&42��viV^��JK�]�L��'��L剚t�n� /t���[l����_�C5��B�Z�kH�DX�!��6�R��𳏌a��w:oT���j��K
E�?%�GcQ�;��b�U��( �Z�N��ҽ�I�"�,fipà��w�B���
^��Ѽl��K��lhi�/�%�24`A-�~k�-V��(�Y����#���u;H6����#=+z��׽Ĵ���F����v�ʝ�}�f��+����3��$�k�ܒٖ��OFL\H���ڠ١qh�,��Ia�\�(l-4;S#��rH���p �O�4#z�+��X����-�b?�5$I���1�4چ�����l��{��ƽ���?a�%%�G�&���b3=2O2z�����斥� �ட��/{��.�H�������%m�݌��?�����neXd��m�����:\��������ף{Ş�5��KK��]hi�"��	�s൹UH(^�h[�!���sAQ�{�2)אO{`�C��5�%��de�vX�Q.2���o�[f����������3�)UL;��+������q�����gbѱ���z��@6(X�&��CY�Fnʅh	�'�����M�Y٧���eNr�ߛӢu��)���L���o~�-��t��{&
ym��_��%J�E��at�<�|_N�L%�V^�@�aj�RC�C#���9�>'�^������q�kOXu���w(��.͙�R��M
ؓ׈i,�"�ϧ�L�p0y19b��}z"�����B�'U���@0�P�'��jѱ?Xs�6f/sfYbu8R�	c�86C�3RJ�3��񳓗�z�K�����b�fL���-p�ߐ2�1���Wu��ᝄ ��\j ���j�:Ji�kS�=E�,Ե��B�s�t2\�<��$�z��Yrb>���tA�/�f<���ɻ
���d��e���!�g��(MfAZ��?M���Qc�TzL��{���Ʃ&��!$�^��22όם���(��5!���[�Q�qV�|��?h���Ǌ�L�ȣ�w7��d�L~1u�(�-�Չ���aU��M�a� L�Թ6X�}b�;~=pvs5���z��k*�-/ � \���=� ��r�>�C�e�z�/eLu?i��p�_Z!���_Ԟ�|�(@OpX+8p7�#?6���~�Î5�nL�	�B96w�X��#��P�S0��JE*��P��+M��4�5:=��gbd�N��,mZ�+�Y�,��7�n��'����&V�s"���;���3�Z�C�����J��6�O�X����x�r�X�Ԇ�"C�q����;������
m섑d!�L����c5�H��+?`@:��*�uN�Y�W�K8�{n���00�BS�Z� -F�L��Ac�%Ә$�H��Ҽ��-�1���v.���<������ E7��D/roޗ̩�ۜ�m(��(+5�),=�S-=#+0x��6���ܼM'�u?�7��u��;���G���i�#�Q���}���?`�(L���~�bj�����2i��b��ϼ=i��M�.Y�>E���l���5�b����9�VIҳ7a��%ۖF�&�������|M��.��*6��z�q�P��C
h�z'�o��Ic��<H��w�6+@�߀��@���p�
@m���n�T*��çt�A�����aB���m� �WSVv~�U%z�ʻ8��$�c6 ����4��?�a�,ƪ��ǒZ�O�J���������]6D�GU�L�o3+t��	��|r�@W�Q%"� ��`'��F���u�L�pm��*>� ���p�����e��7�F%$K��
_X)�<�1���|j�����%�A�=E��@�y1 ��	��~\�(���ڣ�R�����6���r�X��Y��t+�.@��c��f?���h�n�i����L|�v�D�U^=�u���a(���%&�P����R/��l�,2$��"�w��Ņs���#G7�`�`�Q�g��O�2}�I�l�<�^A���{�����ե��!F�ٚ��=O�'�bQh���$qh�)�C;�sV2c�����l� �E	l��0[��������R���W�5�,B܇5����|d�����-+F���l><��Ց�6�,�
N��oX)ʚ�ݔ�wȯG�R�Ԅ|�?�Ӝ5f������g�A����,sTf��4+d�8A����':;�����}�*R}թ�\Ԡ#��ks��-8��}���u����/��?tt[jw����ZD���#�R47�UA}��括4�.��~1x^y	�xN���[��T w]!*<��:9�;,�Y�����?+G.6�+���� ���*��(I��;j�8�^U ����;��pA{��SN@Ng4WBe���٘�h�P���m-Ȩ���>�!8��6���"��3GƿË�r��v=+x++�?RGj�p�!���U��B���m �g�tP]U�@Z>��H�
þkƵ�g����^3��rJ�4�-�����\�Y�Q�4�A�
�}����x֍䙂�ڦ`�3Z�/6����/r@ã�ר��0��m�����\��2Rx�O�K�<�5?��Щ�|Ʀ���|nL��8t�V�0��;�&�E*�|�Q,�)I	*e��>Bȣ!	T�k|�8��t�ݘ�� ��oY��ڰ��M��J����F׃�:�*Cm����gBԪxc���7��'����%t�F�菄j�6�+����I���+�cx��FܗQ������_�x��2^�i�S�,�}3�l�_�Վ���"0��j�BҐ�fz�wN�L���q�����y��Q4RT4MV�S`��rr��(D�aľ�Ut+���A]��?���˼Eưc%��if>���tsB滌/޹�I��#P��EW��K1ȓ)�)9�aX�p��U*�xu�����.kͤ�B�pu(O�x��a����<w�M�CSbBd�pGP{0G�����e<�)镲|�.�wM;i�:�o��+i*O|b�.�	���$��Lm����[Y9OQ��Ǿ1�o�G;c
$�9�T��%��jJ�� v�-񕯦��T��w���~�?	+l�l�-�y�I<�bs~�4r�M�����T�}j(�T��>��؂H�����ft�C��Ì.v�y�C墓͆Z�|��模�zu�0��n�l������>y9/���"�x>-}�ĥ��$.�w/�=XV�n(�x���-��b��G4�xz�e�#���&�]�Hz2p[D�\�?��z�/o��뼊h�T�=PN��TW��{C�����^�u�Hc����~v�y)�"�W@��NІͤ����s�������>ͪ��w���y��$��B���(i�n����$�p�ei��+����p�!�N	���<�i���A�]���2�ݴS��>6Z�������G'.AY�<�V���H����� z��J����/����v�!m*��y�A���\�]p)��
*��iuj|n5h$X/a��U�F=<��=���Y�4nt�<x��+y>A�,��Yr�=�,-�-�~Xf��T�w��ݡwH�7A�6E�d$�����0 F	���;���I+�~��t�ɮ!'�+�k��_x������z���ng[wĖd�?��zb� �V?��L.�9�9zU���ܙC� �$��{e�?�����ɝv9���|$>�c�.!�=g���������6��-����#�"
��u`ܜ�.ݤ��7<i�7x���t�?1���*��ԃx�� e��W�*t�ˬs�s}� A�ѣV"̜�<�P j3�P�u6����R}Çb�7�m�|��������}��W�KB���a{y.��Ĵ��9��RM#i:��+Im�����Ԗ8����̼:�6���V@��'AV>��+���x��A.�N�\�!�}�ȎHغRv���c�ht�,�1�� 	��e��"���X����"z��Ս>5�2�A,'���?���!��񠵥���檩6�=��}��VЦy�I���oIj0��b�1,��o�K��$����~f"��Z%�6EW5=��U�'�f�ڰ� 8Dm�v5�L,7�H�݇T�ҏ��x���}-�[a�w@c��o���{o��>7��uUE9�)ھ���J�.&΅�,�Nnϛ^����+Km�n��CD����=�S����,XY"�`�*�$��D�N�������h^q�m�o됯E]�JF&!�Gr����8��>�ф�x�XID�*ز�;�����̓�$�jp�u�Y�9�Rx3b`�kr�e+�`3�\Gl�3�<]���E�G1�	5�HߩZ< |�o���LֈN�6�F���Gl�����$|�F?j��ܪb����km�Ȟ
�L���7�Ն�y3�p̪
5����.Z��G!""7��;�];&;�C|�FA����H2q�k��}�+Ho�n>��~ܳ���C�sx��dl�p�rx0��äQ%�����?���2�O�~S�P#��@g�Y?b�s��Ϩ�м�!��7vym���b
n�$���% w)��J����u%�ToR�5�(���z�}i����9Ѳ`S�O�	Т�&����E��$�A�������a����I�M ,V���-�z|"7i
�H|���	(+'���|#���++JXz+;W��_�>e���4O=R>�=r|�t�4=���:�x�I9e]_Z�@���+~I��*?q+:P&L�Z�k�L|߇+��e���/��h�o珊 |�%P��P��Ρ=�Nϲu���=�/е!��=G�:�t	T �ivO�!�X�[�
���4T0��B���ү�IZ'���yw]炟�8k.��S�!�^@��W��hoZ?�/Me#�dc�޵�#�8|��?�O���^ _`T��# Ɣ�y2�=�;Ѣ�m�%Pl�v�ɩ�勦Yr���"�����ܙ��k�ux�8h����<�g��>�c�V?dg3��)�'mX�8i�|
�tmy�f˂�*���O	{�Ix��
��('x��A\M�凣���Cj�rGp�^]�͛I|���.�i��b����A��dE����� D��脹�"Z��mn���H�BrZ�'1����:8ÏP�2�#�e2���h�g4��g;���V�`a17�J�h?�Q�Gz	w�y;O:���"w��<����v�v����7K8�j�+F�&�W�|%AZ�����}q�ծMEH�Q����/"�����O��a)�}���r���wL�����|^��q����svU<?u�)��\^|"�ө%�0x-��`y�;�.5�,*�����R�t餛���ARN��3c�|H��a͝`����t�T��Ӂ�x6k��◸���5���#ݒ��J.D���%Ud���`���Gs	��ʞ\��O��m���4w6� }QRk���WW|L�e>�յ����x��0�c���t�%���߿br�sB�𿃠���~i�\c}����b��؊��η
��YhY��[U�6%�:T_}l�͑������H}X����7�$q�4ABW*J�����ׁ�*�a�>�A���S./	M%]l���(
�������Ύ8��`�`�ڻ����:� z�?r{����<6�v>2�t���*�F#s�ZG٠��j����\9��t85���h�r���Pd�;1�X�[�g�5	��h���*>12vb���ۭ���u�T�f���T������[R;�����������Գ���N,�"KD}��{���=���t��a�Ǔ7XAo���G�g�ZlǏ�2b]D5�_+@d�[7�b��+���2�c���)3�^��"�Q�RԶ�G�)b�d0�<��m����=��~��&�������
�����^ͭ&�F%L�~�8�R�'k8˹�Iߢh
E^�A�Eӱ�B��p'�^���A�ׯ�@�|����V�%�QSg!� ����s�Pຮ��:�uB�L��?�0��H^P����
�x��Q�8|z1!�ZNM#tK�a��a��{n͎��Y��W�<�Zp�Ș7��S����B.!ۋR�li�(�;�[u���aa��!���@�R�$a�iK�ຍd>���3����1�Љ�ǲ�्���"�(�	?ҋvɢ��UY��)~��&�ڂ����m����������9;� +�����Lݟ��1i/�Y�y��-�&
9��T

a�>�y����T��|=2]�,ٔ츒��d&���Ddh�������7�,ņhM^muӺ�,�t�O����Z`��	�)���M�������}�Kh�#�����"��fp�;)(����h��ݸ��<���<Mi��x�R�a���v49�����@Ǳ�����
�񓁾����	:r*����eIV�A��c�0�b���LO0t�7��x��<��X�"_ !�Be`Bi�T���**�\|t�}��JΠ�1�u0S��d��اP�F41&ϸ�=hn>�,��Oy�n8�QD"+,�$�w��3,'�+���n� �������v���q�%&���@{f�hw�
)%q
8��E��@�� �Lz<�x`�<4S�}�{>��.ɡS1U��
���i(l�7����͟��J53Sny�Qh:���T��4<2�zVM(_�d��݃���7b�l�˗`>s�ҫ�Hw��N�f<h�Q�eT�Y�	~����}|dəfoa�J��:jv��䖮a� 4?��BD�ғ;k��Ru�4%5��{&�:���w��P�x�<Z�dmH�r��3�Ҿ�2�k���+��!oKۆ�ܘ�cJ��Ɣ������*�Mː���A`�
�H9+��{�!>���Q�X�͟�m�x�b�6�T�|�?l'�\������ÈbV�B+���:V�� JM��9��w���O1?�?�mte1��Xg~�ϧ�~q������D���a_���C)��.��6��c�ǩ'8��1�;��)On��:��]Ɵ/�A���M�B��D�ï�r���W㮡��Ɓ}	���&��q��Y`�U��	B��8��V�9����a��~�8gi��=;֯e�V�T�.��~p�~?�h�"CjW�}�ރ���0�r��EH1=�J���Sج���O�JP��g_��~�%@I�t6�����x�A'�=ё��˺V]�&������H����2��M���)G�qNW�J��Ɔ�pIԔU��'��ME=�4�Z.�%s��Uhb����wIN�O�B�����oG~o�p�ǩ\]pt����^�D�ӣ�{qȵ?�444Q3Q��^�
a(�;s��{|D��,:K�8n���� K������2^U�¬}~����š�ٶD�bJ�pna�s�Q�X���䫗���_xo��g�����.3W�������׌�����W�wμ
�YLj�4p^�m��-�4�v�7M��x���=�t
�_�E-w$����ħ	���(��i|�;�
�o�z7G'iY�3q��ߐ ����QN0��⺂6V�k=���q�#dKؐ�����y��EKn��a���V�lz��GUa	)?{�
�h��r�,{ʖ������f#�����D�z�R������ɼ��&i�5.z�4\�F��b�2��s�����Qm��Qv��^��=T �����^��Q����V�
���s����5U$��p���;"R~�����-�y
�a{�E(}�XH$�\�d��<�V#��@��I	�J�Y�ƽd?|���?z������L�/�e��ՅV��d�'>��*#�{�p0 �GrK�թ���(!ٷ�ߞ���ۆK>�Ø��7��ǈ�-��ǈ6/���[%a�0_lV8B��������%����$L�½�ï����nC��Ѥ�/�5eupd������x@X���U&Ѯ%�r�Ox�H� 8�ڛJqm�[9�O.�6����p�tpS(�u�A�Jf^[�ԷN�)��,�Ɠ��q����4��Lbmuk���6 �]~X%���R�gg�-F�;O��}���(�lѿ���*������PaK7*½�z�m�3��Df�mbtZ[0a~�;<z��х��϶�2Qt��^̱ȴ���'�>FB��o������.�b�_.<Yh$�D�gl�_ђe�Wd�����6�+y��y�纴w5<�D?��wI�{U�+�lQ6{��R�8�#.?nyi��O��M	T�ehAP�M�jmQ�i�'*Au�$��]8�9eJ��9��ڍU�V������g�f�(ֲ�˖Qz!��Y�LD�?;J�*ņ��S?8�����v��v����%<7��/m�\i���Qթ��4ۗ-V�;��;~Fg����j�!k�O�"�g�|ݑ�a
*ǻN'����|��G��33�!B�Th&�oj��ǧ����-����o�O9�4CѽW����:*�����1P��{-d3{au'��3@I�U�)����1�/7c�Q{F4[�&��J��c�h�F�9��z�t�@50����)�lK��#G��[�����8-��6mB�����9���` �g≧.�l�����a��تߘF]!|~�����Ή�����U5=�7�j�W����3P�~{R�F�Πsn&�Mr�迆��y.�������֏L0�	� �����#���t�F�*vGW�	�k��/3��@P�/���W�I����W=�;=�"RG\�O��I�G���6�(�v�#�5����:c嬕q8�M`��T֑*�̘�p�Q� W���2���*k��HM�wSeb�A�0Jg�FZ��42�G2�e2�L��kx8���E@��6y�@�	�3�y0��"�Ԧg���|8j�{�����7�,�������Z��3.x:��ᐱ/"\�5���{W�"���s7��ys*�G�;������^:�݈{��=M�C������H̃�bH֘��l�A�l(�]'��$�;��Ԕ��}���_�E�cw��`7R�d�J<�k�	/����L�;Y̵�B������K�RbC�J7�����P,P�2�p
�A)���o�B����	�AS<��\�,��Eo��R��
��u��@gNfBU%�B.�$��Q⸝T�K��V�#(��Egn��Aq+Z�O�?o	�{�y9 ��|Re^u��1y���0�zk�O���5 ��O�[V|��c]7��e&?w������:Q���z"�{��b�9�����磰 ∔J��kO@��������aO��J1t�M�i:�3.K�]��W >���&����y
V���`M`~�Q�^��L�+j��S����+Ik1�a�����9�����Ў�s=�#��jAg�-p@@>��RPB(�x?O?�14}y/�� �0��ۏ�`"J���m.o���EzKW��6����e�6��q�O�:�. ���@h@��&�a!��k���m%Oh`I�ýK�̑��#��w��tę�Q"K���z�E�x(��������ۑf1�s��fF�Ӣ�|*�.&td��H��=�v�m���'��%��L�oc9w7���9�����!BsMԞ�r1W4�/�Q�X_�w;����eQ�����7�K ��NV�d��WXl���'A�i�����x>ݳ�8g���J�&Q>S%H�+���m=c��S���	���O��H?��{@��Z,<��H�����.'���ܱ�Rr ���&�~G0,r����a��*��eL���$spt�㊡��8��:��B�_G��P�V�ىZ��^b7�(��ƃB��ݓzښ�2�QXb6��l��\����8�3�KU�:F	I�OE�oj� �'}�y��!7q�$��~�E�-d�˘��xCUA�������i<ơ��g�8��G�N�Js��z��E��♉Iq0��+c�]� Ϋ'��1%�b��\FG9�$��N�禧����p���|����eM<F�m"��&;��\�;�dx?��}�g����tV?/?�ٵ��k�+ �yp������������ �Z5y�K��\�@"��R�2�h* ��eR��B/̫Ԇ�O�>�I�Gg]��=aQh���R����*�}OL���9
�"7O~��Y~gӥ�A���b�k5O�.�p/z(�F�h޷�l�P�.��ߪ��k�~�2�j���/�k/#�	��V��%a�v�@����V���6��T�8����������z�w�k�����s����1��QJ��LD�) %��^�C�`G�/9=g�Z����&3�3~k@���9���4ل[<({�m�\��u�K=��B�N�b�%/J�3��%o�#�O�7s���|bqpn���ﳸW\�P}3���u���`�\��Bz}�j�U|Fj|����9Jm��d���pk��5���Xx�u��[HB=���`bفFy����P|8�;�.y�v��:�MU�p7Ož<Z(#NzՀ>3[Ȕ�v;1x �ڨ�"��nǫ]���=Q������#���LqC�띷B����J"̫gE9U��!w��ue�3�������&� � L=
�.àw��qF�mt����q�[�p���xˁ?����F��Ԣ�0�����UG��}�]K�@�+r��õ����߅L�()��bE��*��X]*��ؑ���[M�.�5H��B�͞��]�����Hp}B	0h�]�+�@�R@��զ
�eb�\�˶7��	mi�V��&�G���\�U������4�5���1#�;�tǆw˞~򹊖��o�[�<tT��[Y���.�3cb��+�7�T�Y�L0��r�r�OH��6�:�-��!�'�0�2� �Qн�)��������l_�Ϸ8t�q"�r�0�ߣ�����S�Nʍ^��'��	��2D�`�~;\>����3�c�3�@�{5�����A!Q�m�v�)��|&QH4�� �DI�Mt�r��{}g��Tș���N�j�j	�q�D�8}	N�����˼8r_�@�d/�&�\�8��RfZ~���8xEGF�!?�_N�{ x�,{WBx�0�{�И��lKK��mk�҈�+����mA�>@�p2��
+�b�i9�/J~Liv����Tcj;|��<�p��b:��a͹�� )H��"/24�_���:<^��!sT��V����MIw܃ �5��Fu#d 
+�S5LOg٪��]��q*�V�aY�\좖��$=��w�߽=:,ol����V�+�w��|�h0��Jή���F@��`�T�w�;��~:�ˁ�_�1�9X���2�KT�o�� q���q9\���!�C={_(PF�RR��>P��r@��*`<�0��K�+�̓�?BSs�-�XzG�u$�#R'�+ٛv5Z��]nƗh�csD�b�?9�v&!=���=�=���F��1*@�y00I�,.i������|1nzQ�㗛\�5.hbs({����lo����:�I?S��f5H���J](aW��Zte0�,1�0�ùy��Q+�s�E�QP���kNG~C�+��$7_�oa& "���[H�
�Κ�}�ї�<3w���8.|��p�`�,c��z�n�zd��#�'zv�I ��<>w "�� �=�?�3��#�F~U�y�T�ĕ䨣�$�&yE�ՉZ3K���Ku3�Q)�fU�}F�)�t?��Lt�<z�Qs����g�cS928p�f��aK�����3�s]�pT��M�G���#�)�ȸ�����BK?���Z07�pQ�v�=E�]}�ތ����I��w���R�&\e���L��т2�[�5v�I�@�vV��ʾ������=DT�~Dr�S��Vd*H((��w����b��B_���J-lo�Eh�t|�I�uʁ��omN/���G�"�����
�*M^�qRo�S�D��]�#�-�b!l���Q$Ao���zzܽ�����-�:���� �+���&lwp�~�.,=�V����3�x|��)ֈ��g���2��:YK��&ܶ��|��~�1/���g�w��TN�8�\/FБ=h� 3�Ł�I|T�5<�
�6�;VR)��f~�?z�XN�+�
Ϛ�^�P_+KT��j��c�H�xVr�v�l�C'+�ӔǍZr��=�E�� �z��A��չ��Z�d�m.�2�_{�i�-W�@���𜐒�=R�G��	��Z A�QVp��z����i���5c�Z8jl���{�w�Ѕ��̦@u��~W��|k�ۈ�d+�E,&�i��J�(�ّ��R��E��[�l��_20kr�>&j�V�N������P;;k��c�IW+�
yfGV����A�����d�-m���� :��O�Cؐ�0$��r��@�/��'�a��Mi��t.&;���.���W���Ǜ8$	n�FIp㨅uw�#9��N���Kn�#�0	����9�F���8�RtM?���o+�Į@ij*���`�`M?��ȫ&0�9'�I7��h:8f��M��0��[��:�r��Ft5��j��GEOY*M�~��V�<Y��̲"{bj�H�1��6C65��Yѷ��D�Y���OjSA�p v"��S/�%�Yz-E�G���xkq���3�ɉ�H�%H1_���>d����Zt�z��&c��?4��5��-��M^ΰ·M�E�d��\D��S�c���p��E��}�\3�����e��^�������M�}����%um��R���1�֘E�^�^N|��Fnr_r��_߻��jZ	��1�\�JH���h����r���c� m�#�F!�}:��j�k�'O��:��tI� />�*uzO��fǢ�_G�����yo��m+iQ8 ȫ����]�}�/e��2�����k�@խ:TQYx1��������ъ�e�2�d9CQ��@��^���w��?ఘ����7� 62X)wѱ�6th�+� �ɖ��m����B;�i�X
8��F�>^�J��/j=ƞ�ȃ��'�-LU2��-1���BanU�~�.�J5Q�i�'>��iAٯ���������@�D ���m�CѬ�R�Kң}���#�<7�譌s3	�X
ܲ��խ���vc>��������X�i��œw5�̝��"}ͷ���5"Ӯu)!��C@d��}mIʬ"	Fi��X��ޞ�6��2�Xc�X�[B���fC�=H����ƚH� ��Ǧ����!������y��K���g�^M\DhJ�#����B���*S���}ѡ,��[9�p��H1�upӸ
�ɂ�L���u�v��$	M�2>�7���6�$J�C��W�(�t��"��:V������I�ԮXud�׀�9i�q��-��-D2-~fkS��ᘇo�+R���)�})mR=��\�N7��i��\`|�}�2�hg��!l ԓ���pUu���<E����\-�s�����S ��:J@R�W�����9��*1R,ߤ0J�"B�����PI�B��aj�R��W'V{���A�X�ʶ5�t�JSn��H�Vhw͑([}w͏5(���m�l@H���9E5T;9�DX��ۨ�Q��-Ƞ;�FN1Ĥ�x\8�guc<��0+%[��D��\�X<Hn�dǛgB����}�<���'�t�j�w,��^<��u�I?�<x��a�zq�Pq���Ȣq��E���]�_�<ڤ��❟�^�j�8=��鳇���A��?�;���|���$�R����B&L��ޔ#� q�HI�	Y���Y2@c4� 5�.���<����ɀ;<����\봼�Z��/%X'�z�8U�m�WB�4)H{����	���" T���U}0Lxk��՜[��O�����YQ����C�{��7�G�~-|&m\H�χQ��Up��w�!�E��O������e��&��g �UaTn�A��)�fQ�Q+���K���!9d��8�ॸ*׆A��7����WB�Aa�1��s\�>g�G)g�R4�����]B��Q�e����	�x��46���A�*��k�;T�����'e^U��U�w=����&��mz�
Dg�����_Lj�qHJ��B�1�x��%�y��"u��L�-��g�lᄴ��%�6HX����m�q|�2��:!7_��\��_��@��/��4�'�V�����p=9-x�y
E�Y��Sf匄����:l|��&��]���Z�5���1��P�ᮚ�W� ˅ok ���}%,!�e{�����փ*2E��y�^�1�}�&f��NF:�/J��\��Z�p(̣�MMgsԷ��V`h����틚��9��`�)p�t̒9�ḣ�L�v��U!H���R���]�C�E.n#�̇_%+�e��}ط����>iziVH����8�6Ef����ভ�_���[���A�������a�)���ߜbBo�d�	���4��:�i������Tb$����b	q�B��.(hdKdw��j073��;NWkhc�Пq����d�1����x��0[h�%��Z�t�c�E���Fb/�W�L�U��|o���sm˱7�#`pP�c�~�F�(�+"�H�6��Qh&E��&.�b�A���u���Y�o���Rb�:*��.�����l�35��A`�R#o�r�&�[�_�ZGV�ִ�<Ѡ�H~s/DVbU�: qE��=M���rXp�����+N��1�Hp�F7ңc�&���11�������� ��\��%<��i�l�\�LZ�)i�[1Y�n���2�1�����ud�g��1N��{�a�5� @&���܎��T��ȣ`"���6%a8A����"�B0��sP���8:w� �mym�_�'�TL���xd�J��8]��V�f.6����є%B��6���'Q����|��_���,�4d��s,��Ν�E(��`8�m�ݧ�=!��*���9Ǵ�y�J�E2M��I��6��Pt���c�A�@��[7�ߒ�N;F¹�?2*YW
]JI�袘���فjm��:[YO}����xZR.e�$��WG���0;�Vvk#�a���9_�!툘�M�A���(�VЮ���J��&?� �W^�^�A�raj)Ukjt���a:��iPFo"�蓂]�Xn藀��ؖB&� J�j6$��a�D���$K��xD3\_�(����ڇn��d������Ll����9us����3��X�a#[�Iw�����۵����|Ѻy��]�lb��Sڌ��0�����ԮK]������y.�	�c���� ͵�����͛t� 7�/��|[]YL8����2�o�*��O�PS���ꔷ�q,�P�Z!Pd4x�iFڅ.� ��X[�*4�1�p�����׎�;�����ӝo����D�� �N���]C��]#3���M��A*�2���0��}2@Y�#�N6[�1��+]��
Me�J�Y�@_�v���bZ��a �����:�)�*ʪ\5	����>�����յ 5��S`���QT:�wb�zz����.������������m�u^g.��I�<#P$��ut�)��W4�#+Yh�{�c.O)�J��dn��.C7(��d�Ö\;XдE9�O�|�Q3�`�9��{h��s��o�����i�:T��XA$�J-��/����G��I����׳w*�Ն�m�iL��;}oU4<�0��%d_����bR7��w�(l9�}M�N�<�(�g��l��{'�]=�7o��4I���x^��=R�fq��B��6(1/�d�� \G���)��d5�H �0TY&��.,g�H��v�Fr��S%E���͡��B �q&����]�h���ZJ��B�y�#��5�C�~-Ϩ���褈N]���Y��|s-�8��(����؄�W�;�7�`4�Ɂ�3Q"p��B)���X�3)��k}Tj�8�i[����}��D�Ժ"�.�H�Jm��p\���x�Yރ �_�&�V���X�+= �O���{�l�z���׀��%W��j�yD�^��<�M���p��!/?��8�@F�����dӐ��H/|�0�+qiwk�;��(���$/o��	aT-���`{� ��u��]v�.\\4��e�!G��0(���PdWAfY�b�4������[�S�*Y�46Ggv6����;zjqAxѮ��o��'�k��� iZ����A�����b�)u�yx���|���A��5��=]U<D|D����:ǽy�ݚ� ��Pvjh`��0�ȻB�]_���P�]"������5�ݘ`2],�u��m��Y���x�weR��f�*�����=�݁�^�U�ިOs	�=��D�+;	~�%��:�鍡蔘ʦ�'J��&�l�5�]��P߀�@x�X���2����n�J�Ws��*.�1viw/Y&�w������Q�O{v �/р��R�3^�=��������A̪#�8Dܸ��샯 ��� ᱅q���51oN+b@�H�>�,dH ��6y�#V��t�e���\�Mw�����Y���@����u{���~w���f�}��揮�;������O>+�h~�rϭ���Cua������it�Fà	'�s�2��UմF�dJ�oN27k/Pq� �d���Y5���Nw����z-�I'�`p�$)2e���A?���>�����R�`Մ��,�@-��-�H˰���.�y�j���<�,��6�J���Ҙ-�*o�2w����19LԓBͫNLK��bAU�>m��3a7�I�#եx鐯�)��d�ߤU��x�C~k���C�}��Z�x��։m�~w�>����Cg��4��x��H'(-�)C��*��M(��j��D���|veT�SEt,��r��/E\�'XG�:��(?�!g�ӛ�(�yҋ��+��xC�9G�U��&oz"ڊ7�'|��vT;x�����	��^��%�OV|c|㦤��]��k�=�ڧ D���}�(��5��RD����bO�Vg�UU��;3r���,���~8�-���5��$ /p놶��uȂ����ޞ��qL���{��
�l���$y
��+�u�&'N\��&��7g��3�*���Ҙt���jz�+��Xb�q���m�#��K����Omp��c�86�SL�Wlnt��q�aj7�cVz���9�6phł��X�5�_J���R�` ��5i����w/���6�C���\]��4�-��to�Q.�`��Xu٤1!������<��d�1�w����:���}d���T�،���a%/���ݧSe� �z�{�B���<ȜMp`O�uWf¼
�u�4b�'�5XF�T�Joz�2hL�Hym��n׶$��(�-=�Lג ߠ�OA����wǨ[�����I'X>~�xiN{N�.��|.���P����5�V���KrR�)1ZY���2$3���蛎�{��=��#}���7Zl��quAQw5X��9HA�N }ړD�U���eik�hzz�O��¢ZB�3B��S $�)K������� �O��MC�sA�
��-u�Ϸͱ�n�`�8R��\�*�W����-4�Э3	~�/�IUH�*�﷔ǰ�֨5�4�tY���w����,\�B�?�bb�[����gj� 8n���Ԫ6�*��쇻���j~C^ƥ��OkՄBd5#�R+)�����P�����Y%t�k��l�9�o�'���F[��>�10v���NJX��ܲ��p���w3y�� ��rwo��h������}/�ݭ�vq�l|�:w><Í��<c
"+FQk1M��I	���A�[9��Y��0V�Kc�ޠ�����1�=i��u�VX�q��W�Z�x��}E���氐3Є��c"�:~��Ԛ)/���3��%�Mӌw#�i�f���#���E�Ԡ�7a�Jc�Tf�2,�ݧ8��w"��]jN��LF�:�m���I��\Tce� <��v�}4�ϭV�.�O @�7v��`�PP�=����n���X�����fd�X2�cJ��԰�*.$���#���SA��n<:��Ԭ1үx���$�MCb��p�E*i�4i����Ag�9�ʜ{�w!/FǛ�R��RR�������&�|[7k�p����U�I��\xӣh���ARs��O�B���/�-�G�2l�^a�D_�)���_�d�%�Ѓy�K�sw��C�5`ǯ9����#ڐq~oBw��_����5����R���e��v�/<��1{	��C�,�>w�m�ٓmw�qm�O�SN�ρ8�j�"�ӄVI��Ѣ��o;	��q�� H����6������a���
7d��PZ=�/�)��s��X���.���/����W��F@�����vݓZ��q������iW�k�vR7?ݡ+��x�T���m���D����%��*NC\"����e�����^���FPm��<�FU���UR"�L��;b{̱=�PR��p�X	�u�w�00$����.Ə!�o�~��G};DΘ�	��ZRp�T�w�_��iE�x}��N*d���$��uG��� �fݦ7�b���m�^{Ia�~��:�H6fL��%��}����z�;�"�aq�_&�,�0��s%ف�&�bO�n��9t�Ɩ��SHPu���.^� �>Hk�j<��:�,�e'1�Y0�[غm�s�\Pe2�R����� vH0V�7L���v���ïQ�.)�[��Ȁ�da�Y����V�s�㥩>���J2̣�9��O=v�R���iH�4bp��|	d�=G��#|�\�q�$I������5ԝ;�x*:�ό��m�������w�j�k�d!�0�1����l�.��k�ø�)�H��!���X�p̍ɦ���Ug�|3I���o�?d��O)l/�$cb�1׻�z>5U���Ӯ�OD�s{Q_�m�
Gw�`fuW�ބ W�*�)�ε�oĪ�8�Xn3{̈�����yD9ȑ�2���o�;�Q%r2�}�W��v*|���	ˮx�1 <M�m�@����L#��ӹrj��ש�l9�2�F��m��/�<m���`���P�U�4K6O'D:n2^Dn6��>u��Q'�WO��:��=@I�e5}�%G��ɭڷ�_�P�S���VC>���b �_ٲ�0�d3�JzEu��%���{�����W5�6/��7�,ۖ��Nc� ��o]'�ɡ@I"Ǡ���h��ab��A9`<�('�Oe��A˧���D��Mj���^f��j-�r�`�x7:8�����@v����Q��n���0��~�+�~� 	���K���YG�)���>PeZ��6�3�Q�9�����'!L{���xc������N;���dKZ�,"�Q[;QI�ڌf�8�����U>���0�^G� [����] �|�"H0����pػ�<`m̡/��:��^�Pn)�����Xf��ԡ�ǂ9IHq>]�~[�� ��Edjuf�E�{��"��0�K�1�����Եڑa�SǢ��gL���G��Ҩ1l��E�#i1��J����h�	mt�Bi��ȚD�����v��hj>{�0�F�>?���n�%%�S�!i�v�9k�
�1P������jz|ӭD�y�-.m���N�\F��w���و����LC���T���ej]��^D�i�6�7jK�dY*�Y��d �
OP�Q?_o�}suytw�<��1�����~�]1�C��_�Kw1J��C�QN�Ffݪ��C�0P���s�Z�@<g��l���2P%�^�3���7n����9����$�Įx�5L�l�JlZ��,���"���m\[���^�Gj�>��HX
96�ed�\�c`	4�a	���|��qۙI�,�O`������n&���:.����	n�}��4�;���l����Yr�*c�E�
v��4e�������k� �1z2J������9*	w�yNھ(��nܳ�|b�>���j��ls��!i^nW[@���mo~�("R�4�Q@����)��?O����;���oڽ~���N���~��-a��8C)J���x�^���B)�T��s(E����6�h� ��#���͇�&���fX�up�y��u��nĤ����e�%W&��D��D]P�Ds�K�6\$it.�Hm�U'��3Uq���� Ǵ�˪0n�_v��j��H��?D�켇��%c���LJͿ>�{����'��rL���������&���x+Ľn� ���z.�I�{�w����8(��N���D0�|M�4�~b<�R9,����kj2��3���x����\�h8�cAWs5��i�h�wm�7�+� 6�.���1}r�c�F�Z�[�l�V�K�ԤG&mvi��%������w�����ZaӔ����^7;�~O�j)4"T�=��	���(�1�e���|��sU��'��.�(�DG_�vG��0<v����/V�PEbg�＀�6�K��4<�x�D%l+@V=н�x��}C�J`�f���{���~��ۭ����a��A���Pc�j����/|�R��v2Y��_���J�*5�ԇ�����*~��)#{��sɎ
�ȕ�q��9'��� e�ڨ��͠�?�˭��SpRџF��jFOp�}JV����u��+:xY}�d����g�=��oT��7��4yp�̍�i�>[}��B��XX�����T%�?02i�e"�0����1!�K�.�Omf/ʎ��rNۦ/r�, ׳��y���?��	�iQ��Ds4�롄�ƻ�H,V��*�[�q8��6|̒tץ"�����I�x��91�T��Bщ�d�mS�+�E�W�L�e�X/��l�{h�^-tݓ�g��V�x������Ʊ�@Y���F(
�.q��b�)�d�5�R�B�!j��֚�r�O>��^�u����2}��GNݥX�0�1	�^;D�:|��q�yw�� �C"�B,j��x:0��5{�;�E5�R�6���-��~�����3U;N�UQ��Z�N|L0C������e���?M�.�bi�~��e#�h�>��M��� �_��f1���F����j��=��H�'��Tu��Xm���P>B3{N/��6�N���V{6��c�r�Q(���ƃ�?��*��J�b��=�J��=#�O�o$�j�W8��2�:y*Q=�O�jQm�$�iÐɎWO�ƴ4�4q��z���Mub�1�u|�%�k16u����(�Q]wk�*)�q���8����m�}�M���c�uB`�$�M�d���D��H�f�� KD	��$�{.څ|IB~�p����	�6">�j��HE�L/�q0�[R&͛3v��w�)��G�V�����ڤpv�'����imf�]��� �j�u�x���eM#D�r���XΠ���C<5�{}Q�Gh����N��������@��H]aIMU{��ٙ�0�`2X���Z J����K�ߊ�;���j��(�Eiu�=yS����"&b��V��E��3J������H��/��,\jCj�>����z��*���g����_}	�E9J�=3w�d�܁�f
�8N5^z����e�bnW�t�����UOt˄v��mb9����x!{��$ִֶ�w�����f�^sJa~%jc���r*�i����b%��w�����JD;)�F3*�<�=J�M��oOL��th����´��l/�1M�9u���r*D�w��LBĺ,���?q��������� ��.���j�?	���/ �L�YW}����$.q'r.1�� 諸�F��YŪpT?�t�#���_-�99w��h�*�$4hy��[�qO5�z�Ǥ,�TY�g. E���z3_²�O-@@� mvYҔ�&��c�|��/yw��"}�hU?�61<��� ���~�DM�¨)H3Ѳ�I��ű(H�zk���`~�Pm�j?�x�m�����^�xz]�Zy)#ˁ�r���֜�hY������!�è�]�9�_�[i���NÂ� ��9*�����i����d؈���4��p�`D�\�6�q��q��{-��>���8��J���&��)�.���8ǽwot֡<����� !㯈N�|5���1l�}+˚7g���P�J��ҟ�p���W=�[�Δ"ވ97E�4��It�)~R�L>� Gn���#@	o��6�Cw����7����ã��4r6G&SZ����D=ϴ!,�pt��3�~u��/�v��m'6!��ۿ���=��M���;����v]���\Dm���2��7�Kz��C�(|X;��Ko^E��˾���$�1�� [n�<�Z����!#Y�J�G�uB��������XNP��u@!QH��Sꄙ�o�}.�X��ۅz��(�0�(`܁��Bz���;,Fj㧊�V�&��@+?����3߄5�z�1�R�n��p�CJC��}��� ���VF��
��l�|�ʀ�b�$ɀV�n�p�"���*�ҞC1��,6p�LT�-	`r�J��F~L��BvׁƘdFo�$t��P	�^�o�Z�����1X۱��vMֹ��l���/=� �+�g(L��gE�S�`1��A�}�,��!��+�"�d�s�U�!�쐀�ϡ	���.(X\�[:���n�[ +F�UUR��Wv��w�cqK���
�h�,��Q���#�٬�^�hT������?)Y�?������n�T�ol�6���I̇{l_� ý����Ղ+�<N�<'_]�J{b�j�Q#34�:��@I&�q��K�韇���A䃍�>�D��L\�����Γ����}-��7?����s���o�Q�*H�-��x�{��i��s%H��
	Ԉ�Υt��G.�f+2(�$5�))U����S�6�])ˣ�����F�"r��ֆ0�Hϫ(奌�L(��{��ϋ�\Bz���/�G�i���f7E�R��V�^jZ��d`��,�`�dE�b�����J;Hg(ǇH��Ѷ�%�B^���嚽��k��*(��e@���VO��Z�z��^���S)�u��۬�k�{˷p��W�7���@-�f��t4����X����i�Eq3Ӕ}#$����^��W����bǊ��� I���L�{�D~].��v�oA��5e9�4�E#���z=G!^�5�jr
\�Պ���dOs,�A���F9��M�P�_`u"���!\>r�(j,_�������娌UQ{i�M�Jzw�����<4#�70ޔ+$�"���-8�:l:x��,��{�x��5%��n̕���F6�1�D鋽�d۴�*������'X����۵��
c��Q��Ǫ���u/��~+ٞ��h�
�[9(��Lp:צ�(�,?�:�f�\Q�e�Tw�%W>N���^�9bI����n��e�ƥ�����wD�L�y�:7�*f]U���%��F�6Hw�h٫JHқm@m;�?C�����%��]o#@2�F,M:�!�@=M�G��~�.\e��n�ë�#5���\SBK6?_9��.3��jS�I~��`8�h&���V(� �tf[���F��,@�ugQ����6�Ѯ�n��?]�yc~˺|~^
���g|p��k>���-w���i/ރ]�X�0�n�|��-�ӆ�߶P��9�?�X��
\�·G���� ;�l�hyH�#���W�ڄ�DR3^>QNk�y�K-D�~���k�M���y:w�mO'͡Q���14����EP:��uv f��s@f|(#�>ĩ��N�ru*CA�D�8�}el���i�M#�{�3�4�kcK\ωG�w+5�$B�,%���D��|��R�aڷ]v���1d����Fgvw����&���ןS�)�����he�cZ���*v�	a���U�&�=�b��p��<�q@%��*!:�s-j�[	��*�o�XƆK�*�g��=�7�M�b�F`TeP�͍;��'N/o��")�txC˖G�3�F;�5�4AE�������h��7֋E�Ѩ�p��4d>!��G�R�r}����'c�x:�q.��,��� #�!*P^;mf��,�u���{�@�Z_K�H��Rq�}\W�p-`���ʗ�KA1\��f{
�'B�j7q#W?3z@����v�/���
S*�d,�)�ӿ̳Wy֞L��c���9m��u�	j�Ɇ�l����ɂ�{p���r���L�7~�j�$�"��� �8��F>|�m�[���g�)�{'��v������hz����6ț���d:�b,Y���[�m3������!h�iM��"&=^��:����z����.�c�̒�U��o��w-�:7�ºF�ԙ �˳4��V�I�Y.ԛ_i����ep�� ��ڑ~t4t��[$�R��x��~ς�eQ��n�V�T�T.���hb�<�&j��1B���Y|)��/k�SE�����c�^)ȻAP��C�`�ܬoz������f�#0���6[����l�d�e&�|��G����Jd'�/!ީ	�W��t��d]	y����M��"�r��Z5�ٝ���ziU�Zl:�x{{�:nrU�㐝�.oԢ�6]�Ο
�Κ���M��̷��e�Pcc�cP��M{%�z���q���!䰅ށ	�0����Nr����6*��y;Q��_����t��Z任`
m?n|��rt�6T�~E(�&��[ \�-
E����J	 XȰ���=�;0������"�b�"���-���KU��5]h_ѣ����r7y������@$
�b
z��=6{�ݳ�9�g����	�I��>�<�Si>|UͿ�6�o��p�z��'Ms�5�+�^���x6+��k����h��6��L�	�����l|��f>O��E����[d�9��j½9Q�1\��Q�٤�8C$�G3Q���a�*rMFf� �n�\G��hU�iՇz��n	��$l�(:�27��챎��;�Uz�w�[{��p34��um�;�u�!-�0 #��qB�ܣu�Ϩ|�h6�o�p#��:���k��7�`?����D���)a���2���9�3`����I���eWf|���ī���)B(���l�ld�0m��(o���pO��d�K/_�j��Hi��"�_�yM��F�s��k�x7��0>������*m^�*1��Z�:�M\�!��D���rc�ԑ���~���]2���D}=\:����m|�Ey��R�Vă��s_�� e�����Ja�0����5�X�5fk��]�c:�eU��fȫ�Y�ZO:�^���U�S���%��Ei��D�=��B��x�o�*Q��-wPO�Bȓ���3&6��n�8��盖g���#jV��p��pDk&"��g�zt�b�w���S�1�o�
M�e��]�$og��Eڪ��54$[�_�{u��/Ѵ>��i��q��j���p �dK8r�r�������>�;Aa��v:+�i�����M�e&��I2uՂ���nH�:�=�X�^��\2�"J
�b�9袬�V��%�*iΜv 7�"��s��+W�����Ge+|�|��|�a�-��6�(d�5ڊg~��N�s�j��:�U��ML#HZ.Rˎl�HS�Z,�z�^��~��8f���|هՋC�
�S�]�Y*��Z%b�*���OO^#��k�PX�c�_�)�
P�t9\�ҧ"v�^㒾7�6@���,Z����f=��򜑀r�#���Gdp �q� ��!"y|�{�]D�Z/銳'��4י@g��ܲpQ@�/�8� _�����%�r��@C`��6�9*t*'�ܬ|�KQ��#�k���q�Rf4n�]�QȾ�2'���n��^��W� ͥZ�pS!v��CD�-��+No�HQ}��.�WXS]�&|�v>�����=��fzƒ���
Z�s�y@�or�����5� �b���s���\ZwSc�i����~{ݨ��/h���ur��d[���7@sT�$
L��c��8+ж��"dXr^�����Q�/W���>�mPD~�|��_�J�����2#�����W���b��2��\L��=K���k3��4-�~�	��X��0�Wk~����4�+V��P�Ҙ����_�{<�S��~tDBg�E�}s���7�J�`Z�K���6��q~���L��&���'L���\����j�g��߃
!|��W�ރ���Q�o�]�'m�+��\�ݐ
��i�zvX?�m�40��M�ȭf9�j��t �&��M?��{kp�d�P��U�����L�)�W�ܔ=W�>Z�d,[��\��h�ҝa���;1�D�'"kU@e��(7��I"����u����u�� ���.A�ĸ[�P���wX^o^$ 8X��Y��?N61���pak��S���7ډ��CʧY�ܡ�+�K�(6�6�����DV�:i*��&�q��Y�^m �����^�ҫP+Is���~@�K̙�	p6�^v*9�����p8�,:���z ���D襆���vmr��iT=n�'����P@ED��Rjx2��A���t7v�C
��ں>}f�5z�<cg��#����C��
{\؝�,,��c�,΢9��*+���G_�������ϡ����ų�L#~f�/
�Z��ُw}�'�����KN�⼿z1=�\-o�㎿3G)dm`���"E$Of8�?��̋��.3¥.P���8n� ����4�9J8���t�-�^�T����(�U) Y��Ɗ༟eǄV���-p
Vk���)M�Ej��U�_~�$�l��0�Sy:�=ʣ�*�	��Q_U'�1�3�#�\�|S�4=�.���<_�j���G���%��<�c�M�n�6Q-�璏#�I}Hxk�H�~'ɚ����� UGS��z �b~�R��G�B�2=�ZF۱�n~���J�3�+���=� �0�U�M!,��L��a2Ϧ�|�~�'����Z۫��t�|�3尥�L�o�>�ӱF�CzJ�L�c1[v���1l���~C}��1y�v{�4��L��%%X\:ӓG=�Iu�8�gS]b��"-\\޸��$:��ܔߔ"��jT�U�M��m�?�N��-X؍9��m���px�L���s�y���k�+�x�����`0��Ŷ�Ű�ڪ*�ң��V%ĨQ�'�&ң��	i�Z��hZNC}a�$��"�$%U~��`�f�A%:�i���Y,��.��xL�u�{r���8����C�^/�r���@4^U�ʗ�L��zP�߰�W��Et�;&��@���0��3P��.�y�7�6�4)��V��X�)��~V-g<�H����!rν}韗�ģ�π��*#q�(�譭�)��v�� K-Pނ�i��,�HM���e�w�n�dM��/��Ȇ��k��$�h��W���6��Z�8�9ʐF?t��8�ˌ���U���(���W|�w��OkM���Ǵ�5��&`����J)G�L���}�j�9s��b��Ƚ��[�q�n���]J}�ռ�����&�4�f��F�1��è��p6g@��i䎄֯o�6�+�5o�D���QsCt=��/�F�9�&�,��}����Z1?��+R�esb@������dc'�~!�4�'����������}�7�����}��|u)�|��t��8Q����	�덎�Z���C�3@�~���������2�F�}�����\�'�X������#,���ߡ��Ӆ���n�s�Z'����+ϖ�~�it�@�F�5G-O�^QA�<ä�Y�d�t��A.��`L�v�,+��D�Ob��b��(����F��d�u^S�FV�����'�|�S�R�O�n�X���?��V�cR�
���0d|z���"5�kP�Ģ���P�w�����y��t��#� ���%#��s!��ӯ"<�&�)�vh�,M	��q�=�'����^���)x�������V`����� �B�g�'<�He#��Eۘm�l�O�o����q���~6�����y�����ϑ�JoM�ћ�M�:�N�K	N�����gK�*��`u��I�t�Q�x3�hX}��֏�~T�@����q/�5�"��Ly(aKMגe�T ���M�5���2�M��(aS�!f[�*�@���ekD����^@v1�I�=3������L���tN��������w�a�#�e||�9��V��Ba�]�a?K�/�r�C��N�y˵��!�s�,�T�h<�Ũ6�./JmW�/�1Wҕ�<�!ψ��E�]]�?(����F��N�BQ�yH>�"��ҵKO�j��_@rjc�l ��-Uҭ�*��l���t��q;��6O#�9�aYSp�]#0�<�����dٳoFV.bV���v��6�41���'�'��#��	�/
�����~�n��Iv���;k*"�Ӳ�
�'�>�V�Vbْ�j✑ŕ#D=�S���WP�]iH�pb&Ӻ� s#�F�eJm�H�\~�ځM��Qrr�^�V:G��WA)�!�vj�̾�s����>��̥EJ�v) ��-wf��^����^�)M����|�a�7���0��te��s!�����ptv`S@&�r:�l���yD0Q��Rr�{�@�`�/ץi;�%��I�>¢2��8�#H��k>֑�v�gɍ^�7v��:Q������6���b>��	e���Q���J���B���`�W��Of����&6�Ã��2a5M�~��(�;� �nu����Ӭ��X�7�;{�� 5��#��ޮ�@ʊtxM2��� Ȭ��4%�ښ��R'̟����'B���A�S1]?���HB�6AiحhAgo�ImD� ����jCۊ��#Bvf�婃̀�zڑ�t���MG�60I���8C� Z	���P?���U2VNr�x�i��h�ݔ[8�1r�`$��ƖgȮC��(NE��0�T�)�}ʬz�0��yRּ=&�����9\�';X͗�"+�Bº�N8��&�(������[�8!�F����/�T�ꯑ���쎻X��qߖ9�s�f�+Mq�wn�/e�� 	����J�e(W	��gL.%�D+�����đT�\Wu�l�)u��{|�(��>(�#FLMܯ����~v���`0c�P��׷��0������:\=�F��Eano�i���h�1̌�~U2��2�"~����LP��_�)ps&_n���E�B�$W�ʶ��c
rB�}o ?�a̦��r%��w�R2�j��ɾW���	�-rh��4!t^�{���>ut�o��'�Ww��*���E���4�v��\P-�͵4}����t(s���ݗ�g��$�eR��e[�?��zu����-&r��I�� D�U��dݭ��������Lbew����7�ٰ�ߟr'�{���h:���5����'���U5�Zz�,��hf%+Q��F�2��2(m����g�(6�؜5j!���^ޝ�f#habLx�5��n�1�D%q@�.<�����x��]ًB����r���&��E(��T���fn��M���y�".-J�Ƽ���Q�Nڏ��F��s_mA�1[��wӊ���K����.�	�� ��JL��?�����*Ұg��r��-��9�M8P �)��DC�I�u|վ�׻���������b�U�m���+Sxb��?�4MJ$��Ѧc"��eBlY
�7v',kb�9���-�_LP�l���:�T���R�u:!�R��Ӳ0�P���5Fh�:�4Yʎ�%F��e
��-�%3�՚%
褠'�;�#�y��ަ��q9�>۴ӎ�ь&2�/X�a�{�&i��kqpv��ȐZ;����ZH�������6x������A|Q|�C4V���'y�q�`�;O��5�	1��H��FG������ 42��o"3?�q�3�@[�B�7�75�wzp�V~u&���c��y�&ҳɤ�������f j�m#rR�	I�Q��N��Fk8������x�R��Րb����=ٟ���s�ł��D,�>���s6f_����yJ������Eh�Va>k����/�k����� b�sײ��o�;�$�,P����ηq��)��K��m���O�C4�qj(yX�j�,����ػ��!$Y�S���ZF��[S'J�j"}���o�̟�k��ԤTѡǳr_�MC�^@����S�4�K���Y������d� ��\*��$*B�d_N?
l����~����de�7�T`"�P�}�@��>q�^�2�y=nE{��ؚ��_XF^� ?D�Xۈt��n�� �^{�4�-h�w�\�Q���Q���L��T�c��5σ�q�;��V����B �.YP_���ᣓ�׺�|Q���jyz�Q����N���/�R�a)�Bo<����`���="G/����� � ��ժ'���e�VË�`E����	e�ؕ`Y����(�Zͧ5Z"�����\ܛo�7�4�s�.��G�R����IF���""���=��BQ4$ �g��ȵ���=��ol�v$��"c�����4
���۬�!܅��C�k6	P��A�(: gc�T� +�0�m�������1�qy�T�<�Q��)ˤ�F��H�:�i���&E�dr���bE�Hpp�T|uB�a��F� �-@eE?M'�^z��&K��*�|���n4����/�x�Q�Ȟ����=q�VU�)�=�o�&(g_����D��d�U�X�šmMX3
�߅�Z�i|��^@�׼Ϊ4��FW_�c��W�����.���B��5e^�{�Ktej��.��R��G�ߑ7 lf�g��1#�뗕�$(hE�|ɰ�?4����㮎F����7��@Ky_/#�V��`X_�2Ac�n��-�şU�����:*4��n��1R��~���P8�������B�Usp�T|�Pǻ+	��a����Y�vr�4�%B���*}w"�����g�_���K��#V�x�ܠו�-q��Q:Z��ܣtYYЮ5�n�=G'<�`�(آ&K	k�`|�U��lp�Z=�czB�jU
)���T`Ϯ�0�c�S��}�I��Ǫ��UN ����4�*���oV���vП��VzJ7�w��Ijl�0����w[���Y&c7���1Eг��]ƞ�}01fa�ז��eAb�*BwLV'²�+[�!H{�` �&q�| ���7s�D�����d	(Yv���P,@ݿt������m�ԩ��)9T��%�p�� 8���)u\@-���i櫓��TD��y�r'4.S�OgI$��6��">ק[���-Na����ɜn3� 2��ֺ�� ����ƌA�۟��T�Y��-�
�B�y�?
oB����gY�l��#�I�6)Iz��Fޚ�9����B��#�
�^C\���nt�j��+�&αaZ��e�O��=����}#B��`b�h�@�F=?�c�;OT��(#a��#�Z��A����I��c�öl�'�i�����\�]�ܐ.F�H:tU��o��<������Qt��[Hԅ���03�KH�t�k�U��I�3������^x���u��hT�� �;t�[~U�ԶgA����©:u
���i��k���i���{�m��>��v��pMð�V�ˀ�ԨYі�-����zF��x9����aMn���@d��g;V�_���>�@��Q�y{�]C?%��,~���=�.�o4�}���L�Ku�D\&�?�����O�B��"���pXY8�7�tŹ�e:찟�}C�1��ʟ�%�5��-R&I?9Tř���i�.��ҳid��"��ӽ�Z��L78{��{��ޔc4��%[�ivGCē���
�s�߰}N�L��I��<D���YVrO���}ZT���>�.��B7u"�@�n,��#��N�9̘݈�G5�lʔ~i;�E'�W'�ş��h�St����o,�A��2�0�֖i��z
��������ơ�jXn� �C���ø�m7�(ƽ\-�8E 
������|!��Y�(�ʉ��t�� �:d�c����^� �,�*��O�1��=v��A��C�ݪ�l�v���I�zӂ��cדE*1$3+���t�e�|�}�نc����w��ō9��q�M��%'���⃮ހ�Ee���݃h��B�J�*�pA0��&ѭn#���!p����2��	�bYe���4|���Ga�D�Z̻e�Ɖr�O��771�R6���	�Z��ϊS�: ^(�0.NAR��nӭ���3��T�>� �z����L͓b�4�o��y��ר �'����pƔm�LՀ�񿊑:E3{�?�����=*�W$�N��]L,0���V�W��^�1�����0#����[���Oz��: �z�ގo�`�>T���,��1?����te�
4&j8`���^�
~������3�(�|��C:yڿ��u����D�4���z��q���d�V2u3�$]����k��]�TZOHe�q�Z1p�����4�)���x�SQH,a_;}��V<A�| ���C̮����d>��D���z��f���/yJ�ѕ*�c�Kbڎ���L-f��+�E5	�YyZIZ4��E�㫰��ʹ�Jq�0s>�AIz�O0�}���R`^ �ԟm��?��l�; >���Ukj �K���9��T���LU�W��ݶ�5g�l|=U�`�������7�x��cS��ۙ���V���U��q:�.���(-�o	N21���mh��G/т!�t���v�}^�<����Y�������/Y?����.�Ugk�0��#&<`i7q�
�yY�Zy�G���0-���*x,�֫����'�ɮ�I*aa����tV�Il%�6/3�2 �a� �47����g�3\��aH�s�s�2�8Vf�!կ|�d�e�?Y	��p�G��y��Ȍ T���
C�eeBZry�Ήư�xCwk�*K�.S��#���e�u��;d�b
��D�|�up�u��_�R�:)aJ��k�_�6}�S��-"��0aL����na����uU�*Q�#�����0""�/Ī��V<�5��%��"(�Z��%+ZH�k�,u��a�����-�G�1�g�,N�` �O��f���0��P�'G��^Ed��4���[㾵����qP��b�*��8��R���#��'���3pA4������:'�G.Cw ��i0<�r:w7=A���*k�v�+?vY���gf��h0�:d�G�b-JbM�sc�z�?,�qt;ڦ��?�A��T��:��dZA!8i�,y��HX��(uV <��$��d6q�됼X���ؔ���,�-�4��a�<zqde/����o�ڮ ��HyY-P|i��E��]�$�u�L�t����B�2]��D���=p�3��&="�0%��4���a���.JQ��y�M,����G���ǘ%Q�;����Lt`�-������\�)y�	6�¶{�W�e?��,0�֦��t5���� �Ƭ���~�>0���_E�I���\o�׳��{�����؛��R(1l�U��l�"]�Ԕ��bi��^z�bH`�&����uV&���s��?%���9�
���kI����-�
�V�']��U}�ӻF,�׳�1A��`�*�S���b��C����N�`���.݉%RlJU����T�-�d�(`�4��ґ���ʙ��uɊ���U8��9V���0�]��0*�XŲUv���Ȼ��D�O7��d-~<��/��3+7u=��:?}����<���Y���W�o��f��:�2�?�Eߦ>��o�v�ɶ��u>��Z��D.ʚ�ێ�����&'��݃��g=40��g�B�wC��ޟJ�>��A�w6�����P�a$���Dg�\ <tנr)����F跻������?wW�� {
ڤ��o;�&Wy�bI_�����&����@�$dp���gZ(>h�oӸ�d�:� r��it ��
ӭ�1��g|����)��n�Z-��s"vh1��;#}ce1��^��0n�B�F�wN
{~)�/M�xt���ܭf$r�ڎ�2�X��4�#h�G��!R\j�^������c�-�h쯬���	~�7	�
W%A�c���J7�ط��5r���:g���ʢi��*�*������a��`k�(����ve'�ɚ7bw���6d�s�x�[����K��eB�E��8�CNb9���e������`vA6Dp���On^*{�9�;M~����%�xզT߰�l��pT<��ކ\���5����h��0lY���c����-�ǀ}E����t���3,���"���#zjck}h�jD5�Z�#!(LN	o"�F��Y{,�0�U�M�v�c�)� �L�sl2�E� tᴠ�d���[5��,,�e/�4Or�m]{���\�[�t�U��J���Oڴo7)6��ޔ�Q,`z"9�����h�&�y�\�C=#^y\eQ4H/�8~	2�a���{�/�G҃�a+�2H�R$��)P�H �E�MCCi1��ciԜC��M��r��3f��q=F��/�l?��������k�bX_�
��@SƖ��f9#�c�d�k*��A��_q���-]ǡ�У�eTO�˩�*''HV�ɦ2�)�F���Y�juUca�
���,Zo�?�R*c>/�C�*����������|����Ť#��lQZ�������5�#dܔ���s�P@��׳e���)��H_�(P!�'M�b�}M��$�%�d���{0Чc�i�+�-�����ey�Q UWe�MdP���� P����U���X��yS?\ʊp����$cQ�)���#�.�������h�����T_{���/T(@�^��	%�_�#�^��0�����Z��F����{>ŉ��_)C�
=�>�G['��拂�0��E��|��"��Z�;�7��!ۀ�Z �&�\]�[������Q>��q_�L2���p$h:������]��6ԮH��K��5|)m1PױƜjo��Z��<�Άg��oSq��\�z�'xC�9�&�I�ug�;�l󎽧�k$o�B5���G^Hk Z������o�l�WY0�q3���5<E��P"6|��7�/��X?
}
N]��a��M�b<���nY�w]�H�5��$q���ߏ�+�-�^�T`n���#ǑG`p�{¶��ݾ?E�s,�M$�/����(�ض��3v��ao��p��s2c�7�*��L9fs+�=�g�A�`��Y
�� �|���ױ�Hi�ȁ���!{*�� $��G�m�4y^�Av���%Y)�).�b"�x���8�m��>���+��#�����N�9�5�:C��X°0�@/G#�����b�*�=!���8�Pz�����2]I��#j{v�E��P^k�b�)�U�)KYFd���C(�0�����uf���啕�]�#����\it���ix4����d[0��>��x�E�k����u]��E5��;�-��������!�3�C�`�r̊II~^�S�琅�&�F[����A��/Ta]�S@���Ny�	2��w{��w*VӸv'�l��Q��~�EC"�W��s@�.#9���K��`)~W�+�n�>���Gp�4_ϺP�n����0[hupj�ԟ�z·FF���/^f�L�=�ہ&seD�����ۏ:��Ѐ!�y`���!m\anic�9�e�j�%���(�m�~�'x�k6,M	S�ȶ��8	{ʬ�*�eY��&��E%�mG���Or�[?�)���[~�V�����5�x�ONi��	��������T	�^�T��������lX��}o��.a���A[���*�
�8����=�ک5�y��LǏ$f���H��v�8�+��v��
��g�P(rB�}p��Co�E2@Sc�TF���-�7皇!���+�'{���T�|�EL�8��Sō�&���`7s�r)sI����-&Q���廘�f� �#�C ��7D�)�'4m1��^"^ܤ����>.�Z��5�Ϻ�3�N��P�J�?Ze�[�oj�����U�rZ���2�u�;0��U��T��y��$�
!+2_� N�+��U�-���3�&���`d˚��hݕB�ul6溉Y�ܸm��|d7@����E��^�j�YӠU���%��ڹ1N�z�oi�-�-z��r��z~�����T��[��
hD�'���Ň����H��;��:H��L��+����Ӫ�$!3��P���OP{�^ 0A��f��_)�����P<�#�����[#�82M<�/��I���cϋ=Y�`*#�ly�Q��\�g><��"�3��(�v;
8�E�vA�5���?�� ��ԗD��R�
���>�|C��*.҂ l���G�pߵ���vT�<��]����9�Σ>$�>NF��ЦBӢ'�Q��9M���	�M)ILad�6~��ŁU�Eh�&�y�^��X`��T^��o~���m�)�&��e��W4]��Cn0���c��|�I��v�u��@�k �jЖ8j��\sB�z����M�fV�����Ez���lʸ���m����܈YJ.*P??4�Y+ii8�r+�b�������̶4��$�@��a<�
�cӨy����܂�?b��$�G�cS�.Pb�_"��M�ui	�v�iƕ�K2��|w�-'?�R&`�&�ڀZàSӁ�SS(LhK><�E�z�O�u����o��s��8�9���v���C쑥�Uw䠝�0��>i��������6��"9�j�]����;)T
M3_?����Pd��C0��ʽ�]�N�="�l�
@�Vx��(h�4)����!g�wp�@q��A<zi'@Ao���6���9)��L��w�nw�SD.�<
��;9�!Ex-`Ƃ�?O�_�{�珜�U>,]�^e��P�<��FM�	�5Y�7�ऋm��,)ށw㹬9��Don޿���[h����qE����	X���ZV��E\ }*��$?�K��r}T%�=�
S���"\c���T�57R���,��&@M�j�nQbw���w.�G4m?����V��?��5�A���D?�h�qw�#������>��g����^��?���A�<p�[/�@'2.�1�A�yw�Hôs��*�nEWAO��ty�����6/���>w�F����|x�_�'^�����M�l��@>Y�-RM�E���q��AC�;(�JǤ��?�#�W��32s����}����O>�����-]}o�C[��,�¤���-�Y
�*θ�9-_��$�Bp�^�>
;㦥�j�o���w3؈'�p�l4�5N���"jj0�G��
���0�Ny$)�)�J��܄v�6��/��56I��L
m���}�ڛ����@��M
�ջ�I7��ή��}%�s�%�zPgsd	!j�?���ʿ�p��q�Oǲ\y��ok��<`đ�ܩL�^�ښ�a(��G,\pM ���=��A�����Ѽv��J������m���oľW�
��u�x�S�km��q׌�l�mA�͙)\k��1��������8f?I����h�	��R~��&Tf����9:e�2���/o�}:�i*�a�A���f9w��>�V1�/���
mƖB�
HCR�X}�$lӐ���2�Z	�@�}hFͤ�\堢�G��6|{��w��U	��F�k�w�����
Q$�r��4/<���F��S>xe줁-3�\���$Z!O�Z:K����JRu	�	�o�~Z1+x^NU�����;�%5[�9@�s����a�P��Ѣѥ��%��!�$,�E%�1/��s�j.�3���� �fm�Ҕ�����.��P�r࿲m���)VX�1Y#f��D�5�<I��V��/&Y���>M�lԶ��}l��DZ��XM���<QH,D��j�	�Z��?����hy2�R^�f�z��Y�IH���f���FeX�)�D2>�P�؇���ޱA��#��Z~mu���� ��B�z�Xm�=���矀?���ڢ+y`֐P搈�,m�N����Y%����%� �/Q<v�Д=���n���)l��:�������^w=��p0���hm��_q��QE��n���Y�N
]����IV�n*S˔�~����kX����u���aJ=Wbl�I�s8��=z��d�{�W��z)�Ai��RP��l��ao��}ښ��ޜL�'�{��#����(H8���Nq2��{� �vt�-'��"�@�+P���S��h!�dMM�����Q$0�	Ʈ_��s�G�*�6 ��X����؟�����8]�;Zg+.�yy�Z�����:�SJ����y��V\���i�~ -���3�q�DY���h�m�ˎjcQNH��O�����
`i�b��p�ƽ�[qY	=1b��^�Q�q�@���>���kzA!઎s�m��������/J��RB�"	����9��+�u����$5�� xJ�h�P<�u-���1��u'nRz���>M8�	���o�>d�$L�,P=�%m�><C+0����C����=a��p&(�$�[Y��4�؈@ș1=8�bw�&z���4p�@#�s>f�_��S��A���C����}�gHH�W���` Ot}�I�0�q���#�j<��fbu��QM�.Ze��b
 �M�	��F"I��O'W4Q���������)�Nl�F�nce�2�6^{R	�^��z��j������އ&��S�G���9��=*W�Y��رi�~�r7ó�<A�\�ԗC-y�! ���<�j���`��@(`��mg5�\�y�m&�Pl,�,��o�b�1�5�k��y�h����i�B�,S����'J'&��Y�������|�{þ��}�6m��-7�2��[�W�Uc'�,�8�G|��;�N9P�<���6M�ݭ}�f\k���!�7���ϢՐ���Yq���	��I��<=	ER��6u�G&+o�W-�M��2�����kg�ׅ��ɂQ�'T�Xg���{��n�}ʀ�.��!��tcK���W�H�ynB�L�{IЄxJԍU�2����5�%�(���-iݕ�U�?ߵ�Ca�\�1�o;������"א�k=:�Pq\)��܍\1�xݎ��p�����Vi�����㻸�����@V2�{΍�)��_!T������;�H� �׭R􌄻�@xO�c��]���#��sr�OWQ�VmB2
�C
d���<@
�u�Lh�Y�K�*/����!3Ι����T8�ا�xt)�� ���7{{�[����˭�oQ��kzL�/�F��+�=�Q�U��{k9h�b�3ܨ�'�h�΍��s}C��kX+1>��VU�	ihք`6C�p�G�e���V�@M��WBz��EOi�Pt�Ǧ���0���w��G�4j������ɠ��8iw/]��z� �-�i�L��{�Y(|�u{&��� �1�e�ԭ����>9��I��CTyS�#�M$�`��7g9�V�6�ӈ� ۂ*�qw�uR�Be�xO�Ih(t�%'V��� ��H!5��m��HJi�%:Y�آs �v�k�����I?vwR���P
]��왪��e�t������X�^gU#�\���ƬOf�n�q���m<�%"��C�&�6�0x�1`��٬���������sΉ}K��)�)�o(]�9f�Z7��i G�Ko}�Д&P�S��wI�kb>1A,���ň3�#fyQ��y��6,W#��ܫg{��ӜX�D{��y+E�X���o�%n3��8ccFo?^ �gЎbf��"��D���������}/"�`-о2
���O�
<�Z��}\��.���4�7qI$b�--��J��*9�>5x�Q��EI�`ɷ��":F�\� �ĥw�z�et��LU�蹖���3�q�����|_�˶�ʔ�5s�"R� ��Tg�� �E(b:C��AxY����[�?(Qm�Q�!�)\���J��^!�ˬw�Y-��]�E�C�E:��Z$���V���e�����
y�H8]�k�}�y�$��_���=)]���3+�,�ImN�{N�K�J:0���� Pm���P���.�1��$$)�N�{c{<Ew��Ӥ���j����9~�L�w�����?͂z��);|����sX�!O�2K�t��o�i⯐_��T��wo�j_�`KF@"�E�x0W���ln��� �.p���ђ�]|le�۽�+e��*SA�K3�4$P[��T}� ��MEC���EA��$w��Pn�z�J!&�{�?�oRع��ݕ���J��n?�#�Ƞ2%���L"xEb�`}�[u�SE�������BJ��(�Q2g��г�a��G���Kl�����Q������j.���5nO�jO�\��o:�8�X�N��}��j>��ʮ/�5}�i�9�#��	
�d��#��p���x#eF�'��Y؂���ڊ� H�!j.E(h������|�CY��p�W�|����}�	h.�Ž�+[ѹ�K�'|�R=�iK�����%�a<����o	4��s�B(B�jl;(�%2�2�]��R��"r�8QJ[G��ޞ8�'�X�X�?!�����Cc�i����he��\�P��:
S?��6v��u������+=[1�	<w���/.�ìF����*Q�����KV����*�GA녪��n��գ��{ȃ~�r#KG�b)8A��e�B�q�ڬ�+G����#&OG��ƈ� l44莣y��xQJ�`�q d�m\��\*K���l�$��ED��]��2��a�.ƒ�Yˋ�S�;y�[Ugo��;��K��� gi(����(��ݦ���}��I�9�oK�(�R�s�t�×y����	������j��yQyfW���3#��cu�~�F�;p��Z"gF�A��iZ��=rx�+�N����P����S�ݹDY�@���}�,�;yӆf������1j?������6et�H�5|k ׁ�Uj}��|���N�	B���RM��%��Lo����98�"ÿ癱�:�t�.-,"Y�Zy��W�ޘm��4	��į��~3E0!��8����{�x`��k��A�إ��'#���o7�v�8��Pv �2�T8��&�eK��J��(4��2v����۱1�ӱU�	K	uN,����9O�oM���݂ �+6�7i�%k�K�C0�~H�V���'��yR�=4�]k'��&��$#K+j�}o�
A���/�>J(������>aƠ����(o��;9]0r]^n�`��FX�RI�)���q}��u�ʬ$B��7�"�x��d����s¨�=�Q����5���St���^%A�����}̕7 ��?��<l'7�>����;9	%"	BOQ�(_0�طҊ�<&`�$��N�)���%�@9�|�߳y"��,�B��ې�ؽ�G��І)���Q��6:(%�KsV|NG�׮]a�U�O9⼢�?uZ�$�h>ˡ{�56�Y�7ÞZXm@�)vc��{��C4�wfBM%n�;��z�)��4 (5�~k}U��3j����*�@�ƒ�L�E/�G��5��[��H��ME�k@��J+�Ke�\z|���"�ڑ�ڽ�Qݢ:#���s��M����jӳ�R,:���Ň�\>��u��;�`�ף�	�Ϊ!)�$@��³F�"n���Nplř7��g���Zc�ln�{�$AO=lˉ�z�Q�l��rjAc��ĳ\F�o��MV�/Tf��'7��"�#�������˯q�����	[]�����D���͝��Gm��<��o��Bb�'7�rxr�8y�����+�d�m�j�6#L�����N��xQ�� t���I���8o~B��3�g�!Cg����a��.�T�'ms�γ��kN3dhB
�H����,{Xx5w�K�?�NMP{�����iw�Y���� ��'x!i"���<�~m��A)�L�Fh���I�@������gi�ƀ����Dg�ý��T\�������B�Y�1�*��������e�[l�q�x'�Aڇ���>�\P}���@兂c���WZ^a��v���7Ͳ0��[d�g;�3:6S����ǩ�ַl*|~�@�MM��+)�Yog�:������ȉ���u;�������O8��*�.�r�qܯ'!ܱ>�x���LQ�W��o�_��+˕��ɘC�&���'|�N��{���q+Ŗ�Ģ���]`���ʽ3|�so8�d��a;)�U��}�������/� �s�v��m�s�Y�n�e�W���������;$��C��Nx-���yD�G�=�_�8�l�cD��7vǷ6�1�W���w��"��`�Ճy'�������.*���tP�$txZv��Y���+<���=0�g�:vޏF1+��y߾P�X:5�LPg��^���#�q�Ɋi{E�1r���9�gFP�ic<������Ĕ�o���	V��q�s�dZ�n�s�ZR�9��gz�``DJ��U��]9�ZhԫV*�'��זu�Ez�sz$<Z%ψ^|w��T���$��W'ٕ�� �jl�#�`w�NpĬf��ѽ�zA���}�yMCo�0|ro%�2#$3yB����1�"�;�\�ב%?��q�	m�>>�K"��1VU8�X�F�������y�Ϫ���u�s�Ry���c.���!�nN��0������O�q���t����W����@��-<ٺ,��ԲTyF��dy�8��7�Y��M:�&Z��Ct��f�j!��������j<b�v�Ǡ��/�u��"���Yk��'6�W�fžM�����t�_7ݦ~oV��x����Xun��ợIA_Q�}($��""G�'p�V=qr��n��$r"�����l����uGe,i�z�q�O-�5��0�Q��9d�#����4
m�����C�h��8R+���
܈�;M#w���;(�3�,^����{�M���U.���Ղ��2Vj��d��XT _׃--.-�#�p�#��&��I,8�.��Rg��gu�NI��=>Yk�E�2�='����7�����+��/⾟�������zk�n-�ܑ�` ����"Ny�?9�
��>���|p��r~V�J3~UI�b��x"a��0��@��#�).�(F�3����]�v~��O�;�r�8��ӛ�b�W��� nK`ޟx=���R�ؘ6����4{h]�h&@Ԝ~�L�5ő�҆*�j�0�1�M�#0��o�:���ԙs�L�H��U̳���:9J�"�琳{5����%���v�1˽kԣ���	�S�$���{�M�V�0�=��5�{�u����4~B⚶H�0�����t��3N"�ү��p ���$a;�KaȖ�=XGީ*ޡƬ'6�$��n����f����G������웸Da1f�c1=�^j��Y�"|`*W�ρ�8�,���.��D�4�vwR��o�D��/�ף��4A4�W�d��mtX����&Pl�������Jt @�۲�iD�^|{�:�X��ޒ�����2�F^���%�է�4����C����m �4�Ad ��(+u����s�}�H���|�'@6��r�����fl��sF��:7�\�cX�p��$ݔC�� UW:Z߳W���5%9�sBJ�VCit�b���*6����+�e�q1�N����]My�uQ�G��̐tS<��5Z��h�)vq�vS	�~0��Q�:���{�> �<`��M��AB�z�K֯��~Q����ԐqCN�>�T�/<��B�A�k/Sl76�}�4���� �\yDq(m�Ƕ,T���-�����@���F��tR��j����g1�%[ʖ�澎Z)zV}$�|V]W����ۻ�R{���zDǜt�uP����P������)s!d�ҿ*��x�/l�g� Z�q��~�Ͳ��>ԆL��E���=j�)G� �z��K�	[ʦ�&q]���;ͣ�p���hr�-7������~��90YU�+��ϼ���oAo��g������m�8��LU&�����O6h��9�l�v@b�ŧ�
@K���	�:'�k
W�e+�J6D+��4����7'j�AV.�̑��0%6姽�n��(��v~��qB¬�1�<�M=8i����C,ė��g�z�0�^*Gl+�N���F��	��-��Q
���tJ�Ĵ5d���=��7۲59o�h}xA�PH挾�1k��H}�W�a9F�������L��'��7�Ϛ��R��%G��HX��4���?��GT���ϙ�����Ьd������Y�7�hY�v����'7!�FQ#�^MQ��T7R�^��C)�hc<�9�ք�	c;	�}��g���L!�EǕց�%i��z�ܼ����o1t�R��=ܹ_�-ʭ7Y��pE�Fg}� HM9��$��rL��z-*И�ܤ(�v�>�|j9���5b;���rF��.��p�|���UO�����b� q�%�g�|��e���?tX͢4q���po&�=P�&�<�� �;k��Y�7�J=���.��&��x��������m��8���X�N!���;�]�l��r��+!Q�Cr%�C�9�q�:�	�	ZWQ��t�����Ӡ�*�N��Z��RLdEFl��2�y�aK��m�
(S���_�.r���ׯ�R�^,�m�&�d�f�_�|�q��N���� �jp��BE�0���Ϧ��W�2m�cK�x=��Piz�`�t��ځ�I&�4�k��.%:wC���[+���Z��J�M�2,��=����+h-L����O��Zv�kEM�;˾�A��"1��.�Z|�V!8v'$Ei�WB�����(��7#2��J8���\���ͮ��Q9�W�%��U����]@�2��ŵ՟���u`zz`����8�E��B�a6�u��n��t{�/?*�<�^��Zk��Ť5�܃�� ��j�!��x��[?�qVv	of���0�o�C����H8�dy���L@��^��^�^h��Ȼ��E�~ާ��O{!px�X�A�'�텸8C��5O6usU�ͪr���mQD��9�I��_�=����K, ;3��ON8�/�"�spϋ[�h_B[px�3���i=LR+f`>.F��������\$��yVA�_:���[�.��U��A�n)�J�罕��%]���K��t���\�Ѥ-����v� 6<0��q� AI:Y��`�} n �:d�S��Y �z^�y��+ �>��,��(r�﹆#@�$q�"�Ş9O cNY�
�!,X(%�������3@vG�2@���j	+�d�~�A�d�zY˂!�l�O���i��Xs�*��$g%��_��"<=u��;��7)]�,~�ɩ���� c��4��b6�_���#J��H=�O�]�Jd�Q^	�"j���}u2�Sͦ1Ȋ�B��dt8����g����(�Ԫ��b��C徭t�t���
w�޼�/��4꺜�R߇���oA.�	�k)R-��U��0Q��^}ق�r%�6m;m7���� |˩��٪�_�_{oU�W�o}c�S���^���$�� �̑�S
�߱�bE{�l9��˧���w�E���q�^A|����H[g���U�P>!�@ Rq?�{���[�ς>����ҝvzj<��i�~_U`kl��϶����.p�U�� ���:R����-�X�6V�D�O�����Z��Ob~q,��!�Cϲp:�]D���{���;�h-x��e��"���AI�r�M����	E� �Te}��2$@��,:���Z��εv��0���K�M���D�^�>�"�n��@ �gu�`D��y�ld^k�^� �͇��o�o�TW����� �T:�5�vbӦ�����S�z#l�M9mˉs����~>a�T�o,�}�flxju�}Pz�%���WՐ�I���=;��[E�(�LCgZ&<��Vk��i�=���uw�N>ש���n��� �D>U�	���A5��r��Dʦ
���������6(YR�����+�#ݡ��7��^����'`��aF6 �!*�=�BmI}���@v�ӡ.N�j9���d�4Z�,[y�fV�'� Ʒ�+	a��27h��S���Iչ.�ʹ�{�����L�L��S����D����h��q��W�Jg�Wy>��{9u��.��N��`�`ON������vQ����P�Zx`%��p��E�U��:��ۀ��,�𸔂�HF�����A��Q��!��zF&��_N ORi�*��:�iH*qŤ/Y�t!����.�h�o�֧a��+�<U�5�FP6��Y'���x�OQ��	?��o��Nј���l߀�N6 4��;C!�a`���K�~'u��[���ת/��U(8״<Aߑ���-9akʔ���Q�Xv/N;�a�AS	2J���TxX���0��ؐ��ϻb7�O�xoΌ��P�_���~����ے"�lr�"s;��]�DJ�G�
��V�,�<T?y � �m���cj����5Iy	8B��&�� �D �y�/�H���,C&)��!t�a����	�F��s�f���Ava��|�x�8�݄�b��2_6f���"Oa��I�q�� G�a?�����]�Z��u���	ur��'�x6C,�j�w8kd3R�X*�������/V���$4;�5������D!�z5�M"��b�9����$�N�4�p�Y��4E�yh����|���$z�������s�D���'�(���N���Hm���j"��m~�b�?Љ��'��~Z3E�u5c�啳.O"��O��4����m)�������~8��Ԃ�jf�G=��g{F��W��?{�a�����9�_?
������X�p��܈l�{��3q�f���x��ؿ�د7�	I��qB{��?�S]K��T�㖠Z��<��lr�e���1�h����<��ɳDJ�Q���Nv%&pS!�`�e����,��q�"�4۞�����~�2`��e�׵�gOI�ig:ߣ{���~�����@��ߪ�_J*���j5z������7�#4|��-D�D����Is��,~5�]-8��4}��Y-��U�����7���}/)|��[�t�ap��PBc�S!�����|�����Ul|p��?@!�^�'q�.�W�.����G�r��Zk�wr S#������j�1����с7(�n�[�p�ل�ޮb*���S�-j�{�$�`l%��'��Z�Q�����3�SAn��fY��n~�9|����c��(�5ϩ��'J�}e�T����a��@�,�FTvj5^蜎r:R�P_�����c^"��h@�⮁~THs]=�������O���W�xh;z��g(;��Dm[�ho�ɐ�S0�������?��2��Z�Њ�$�IZ�;����p�|���\y����}�?�fQ��uY#���� ��I���.���ye��M�7�oQ�#�,S&>��{�� =.Ɯ��P.�����z�������\�C���W����6�pfF�qۤU��{�S,�����nY �������1#ֻ����~Ed����C�ӣW�"�-�ԭ���#���%�AG���	S�&rX�W6�'��d�\�+�M#��(�k�ցm	�sYw�P�?����l,iYJ:`��z�$�'���Ԏ�U�ӻ�EI���h��4į�Z�m#�S�V���ˬ,C6�b�����2N븄�ϰ�Ip�����-Vo2xZ��I�n��D˪�|��8S ��1��.���G/�570�
j]� yx��eVα�	�ui�f��`�����Yr���Ѓe�t��m=9�ض}�y��4�U ad=��"J���E_&������nr�"�E|��o6�T}����1�@1�ȝ�Σ��""wvS��IEkB%�����Fv�&Kv�F����}��:�C'����c#]���x�~�E�E�t���X���P(�0	j�$EaU�ܦ�,:G�:��%e
tS�gS:D�b�*#���q�z�^��\��v���nKM� �6yA��t�Bu��Y��:h(��*��_�6m]���Ǌ��+6$"�It��f��p;(]yG��,xXV�7��D�6��i���E���h 8揧�2����#�cq��IV�v���Yu�=��h%y��_r�������D��R"����6�} $�̝2?�{�ƍ���x�N 2���&�F6v֩�m��zX/�2Y
ߎ�E�Z~���I�?�+�S1(������=�L�L؊9��6���lҺ�w���,����1xZe��,'/>�!��uaF_Hzeޛk�Q�O�m�n���� �7�b -<̼�M�r(��6�⣁�SX/3m��G�8�)�@l���S_��$����{��{���a��Wk	k$�\羫B�j��Z���ɅCC����Xp�x����ջ`�Ы��M�Hܩ�Z3Ӑ�2Y
pE�S7��3�STD�_	�Uզ�i��9p��ч%� 59}h���4�H��H��u>�hM@�]<<FJ�k��+��J�5�ǋp�U�6ä��N@�~�/��pj�9���j4\��A�7��X�mfI����N,Z`��떷��wsz��9zy?�y<�p��.������k0�B��A0����3lx�E��`�B��u�76��,�~*\��=0��N:�ϯ�/cݪ��N6�%B���gU:cP�X J9=3R��I���*�X4��*Dc��k��ɖ�Ÿ��i���͹��WM����̼ܦ�Oa��-�[����B_���݀m/IN��	��[g�奰�5��mx��2�.��2������b:Є a[���u����4����o�s2�st�WH��>Z���H�ǀ�`�jGX�V?Z�
&e�k��kD�HC�R�V���rI��ֲ'GT��˄T�#�o}��^�Y�*�,s�FLbxll�	���l�3�_�gB���k�P%�$/)XNb��Y𩨪Z-1��T�Ho3��M�.��8�07�c��_�ȧ0�l�/I�b<�y�z4\��B��å%r=>$-�m��Y�q��@�rA�xNqH��jJ8���cY�cmo�B�B�y��8�|��9~Q憎��%uP?Ofȩ�y:��@633F����w�r��C�F���]e1�H��xk*�Bj"�b��-���q����Es��D�K#C�E��(�����?{#$K�T���J"�������h�9���
zxY��P��^F�َ̓=�kGV�����fq���`�A��^N[��t��P�W]��s�1�o�;ʊ��Y�5^����26�~�>V8�H]:Q)5ý�\i��j'x;�}O+ػl�m���֚�
�)�_���V�V������L�k	��K�ɼ(M�6�|�0�?��Ǭ(�"{ƃS#���<����D̗�}���@��dK��3�H�`{�F~/��]dU�|ۡ��c�jO��O�յ��ub��ڻ=�m�Ϯ?��|$��� ��k�&�HQ@?ԷE���z��f��9([��԰�I�{�k�=�З�az�pZ�(,ۑ�E��>���L��vYi�"�<'�2/]d�j9�v�1�<X�":��Y��9�u��^qD춰7۬Pdŧ�I�n�z4w`ߧ�aՌ�lYf�>������{�������;U�1�|�+��If�Ш��o2G��CN�T�Ab�v�^��2d�A[��L�?=�G�0��^*��L��i�`nF'?��F��[O6��ph%��OB%���NU�*.<���R�`̕Oӱ�6
��2%�ͧ�ч���3��#��r��io*CE���9[}�ˋͤ	G�=��*%w�V]a]£�
ք��/daS�S��VE!W������Kf(�i�i1FobW2\���6��d������ T@���^�.�
�$�X��Bcr!�#��������T���UB=�k�r:��/f�ǽ�j��٩{xS��lV�����ne�*�;�J�C\BN��/����O �^�� ~b9�F�u�2�����ʷ��ZR�r^J�K�OZ�����SfFTzD��׃xb���7��}���]t��,�-u������G�4[:}��8J��T�Z����� B�v�A����-��
�1�z�"t�%;1/��!�q�#tW�fp o����Oq�3z̺�}P���-�m���ܙ\b�9�<Ίt�i�
��"��H��.�y.=vc�\aUE&�|2S��������9-0��ÔJL�
)��+���0���� ����'�2�V�������З^�2iF��: ���<a��w�$PCG˺��S��B��H��w*ް����`	��P��:o�
��DR�
�q'�(qe�ZE"�˿���j�|��%�U�Q-�n�%�]q�ݼ�6�ԽU�]+ġ�
���9� z?�}.j^8��"�\�����Ρ���V���yA��ËZH�a�Da}�z�0$V<*y�D�❁��q|ҩ+}"��'�J�9:6���W�� �! D�B�"���C��û<���n�l�VYK���I�ϫ�7E��Q;�(NFέv��I��=g��s�ʀ~z��YݪY8V��fu�q�������"g�'���'�BE���S�\��H�V�@�
��[��_�y��!�Zh;��+v����6aA&��O>A5�rJ�L���s�Z��<�3��3��wC_�f�M� HpO�FN��p��ŵ����jA&���e4�%@w/@��d��a�N\ϐ�ժ��?��!uR��NGз���;el.��gp|!���٦S�c�Q�����q�r������������V�ɷG@�l�-����t{�C��:���Y�u�=���"�D^{֜�����@hs��n�f�B�m���·)�&��3�"z����JC0Ci3���΍�w�w��l�#�|c��%��7/j�Lo��5g@`����'�߾S �ɖ�pn�����O�m�h�.�
$�s�pF6[b�.��%hP>�{ӂ�i4%�8��9�H�eZ�*=��.�T�)�4WU��R?�"���_�����=l��)7��'��K��i� DsԬz���K�m�Tv]?�+m�u.Y��
���
�ϓ�����&���r�@�w��>�4�v)g�~�6衜���a�1��}x������m^ae������"���#�%̾E�<��k�Q(��MH�٘�*�!��)�Ӡҥ+�^~l<����%�Yk^��R	^Q���ӊ�F�(��wRͮSA��@�/��H�\^NkK���H�Di{���=K����7�SM��z�K	��O����^�G,MI1�����%|1:5��&���x���+�XU	YuK~� ��h�ы���h�T��֢`a",�h}�o ��zw!�����݀�=8�I�O�r<	^�?J��+�����D�x��1����D�#|_��	{�m�<�=$��ү��+����U���C�M__?Rݚl���ȓ��.`��DE�7�Q�9]��W"��K]�S���(�ر{J��h3���+�0%�a����%�7ip=�F���y��^!�?c�p[9j��T�����ң��,�_k�U�>�E"�J��a���B�Y���G�I�D�J��+>�a)-������l�B:S��k
[c
O�{��
�4&|x��f�v2�/���-2%�6�f���Jzo�J,�I�mM�0��O}��Ճ�B��{��S���z�f�qaՎM�$���vA�{tbO_\Q�l扢��Aqv�EĨ��uT*�3,���GR�7���T�(OA�������-�v,v�P�!�r$���A
!$f�q��qx����}��6E!��o�p���T�� �c������y�J��	���;j�aQ���A��� �N{R��R�bI�	�����BP�fh��4��.�����ޱ��Vي��5*]�͆cq(�?�ݵwS�Rg'��"�D�>�O��2Y�x��i���~ׁ�Ե����G<5\,>$��\����擢-�e-�M�k��S�@��br�)#7�R���l�� @�R!�'(����By���L���F,����IW�;)���@���^�AȺ���F]�Է ˿*���.�s�}��&�:2	n�1�)~*w�I Њ��.�ec��A�s���r������6�OsA���^�~�W�����q�1KJ���[�F�����q��t	kȴ�-�vy.k\���xh懑�\viRG���*��	X	�X�R���G�a�E�+�E�k�#��q� /����= �!'�����f�y���a��RQ��j���[�Ax�/�5���ŉ��(�g��>�����K����x���q��{
���Ek��s<e(�/��`���;|�n�Պ�6PlO��rȤu�88���XYܿ�dQV�)a��d�`bqJHiZq�	��:�*���s� ����)��4+�cH<�vR���g�R�ٕ-��)xf��E�!��*�����Ǧ�>��  J�]p�k����͈N7h�vP����t��IK8�>�#�u��SL\����~ +�q�� f��-�#,&N-�%^�:CK�}�����f[��V؂S�3Z!��;]�	���0�F����s� HpD���Kɲi�6N\�m�c�F�ǟ�B�u�1ח5�;��O_�~K|��]��c����3L�~�k�b(�V�ޖ,��Ђ.>G���x�M�Y��'!�2Tp��{���|f�w}5$��U6���/�$�����!���K�Hj�W����ߗ��5�6H���,�zΡj`%5�h�,�����Ijz[}n�M�X}ڛ}����"D��N,����8so���*1��+�yK4�����v���"<���_�p�*���ҙEeW=�����c��������x}�t���O���.;<�'���-��(�=+��N�������dϙ�U�4{��a��w�� �Џ� �'���
)�5��G�%�z��s�/����*�oh@k�8�+c^�!T��q6,#x5��d���gA�sỶE*r�^���&��E0�̼�P�+��T���l%�p?."��a�X#A뻺֩�K�yEا���L+j�M�~�xS�_�.���S��{�dT�<��ݡ\��[pz���� �m�q�!a%��y.����F�Ʒ�Gq~3�,��W���ǗZ}b�PT��!5r�{�#�p��
̅�Y���	�G;o���t�?�>6���b�!<��W���~I��cP�O�O��Y�T���F~#&�fb�O31b@����k�wX5�P�o�7+�	��ygذy��j�f�u��)��4w��b���6$[k!��i ��ḷ��`��`kBټ7C@�m����c�7@{����;��'δa��#2��9��	)��ŝ�ٲ�E�]]*|2��A�An2��${+t�ДM�a��kY�zL"����ZO�a��5��GE�f��l���n/��(��핅g�@s���3;uV
��L�<MgM��`.U)�~��a~t:��@����$v*�����'_��X���q�u ����]|���Y�����kr���ml��q葵4m�&T���@ۊ\�8�Fo�=_�T�Vs{H>'�?%k=�n�T��`�k�I%��L�$�- IH�%��SMU�4�GKᯬ8"k,�m=��������OV���Se64�L~��`�UkK����T�˾���4���J��mHR1g�,�?y�t���ƗX�B���Z�߲ �Y�] ).9�͓18�%��8�$ N��߼B�0S�o��1���_�r~&$4^�:ß=ۇ��(�9t�īֿU�����Y�PY�+�|��R4�m}����<:�Po�]�+��
�H�hT[�)��\�y���� ��o����Y�~��nDV��G�5Ȃ
�l�jOi��tA֐u:(V����Ƣ�V�I^J�%��9`F��1_qӧ�?���nvvf��KƁ�}� X��C |,c͚��G$z=��#	�=��-x��?G�q�T��5�KJkK��L�CJ�s� ��7�������9�V��}o"8vI`���N-�Y��B�L"C�g<6��	�)�1]�`�Vm6��K�Ǚ����j��D�n�'���g���6�D?8�����Y:x2�b?����7+P��G�Ȭ��?�T�����Z]�2��/��}��!����.��� �ϕsE�72�<M���L��g�俟���XTwV���ښh�^
����N���єJu��9���,<Ȍ�@̔�\�6T,�^�P�S���
�q-gzh
(��O~¤�B�s��_l/�(RH!b�����Q�삵��Z�QO�?�>'xR��`U��pD=o����#�X�	1������m��U6�6�2��&M�2��#�_k��H1��_j}�z�^��
�.n41��Da��6��e4���st�d��H0��Q��㏡��ek�1|iC�~��&N/=���~����L:���B[t{M��B����0*,D���-*�+��u�o�;]�5А�o�
J~%���p94����s�-n�~ Q?އ��p�����r�D�.�P}�*$�<��^\����vD��nTZ#���kk��؞��3P�ѱ�[�M��'ૄ���an?�p�s2,2α�Zb��ːa�<k�����K8J~�?����H[�e(�����&��+�G$��I��E�CF� �,פ?��0
xmK&Đ�0�/W��D�N"j?х���	"&)���d���tvJ�����ѺTE{67�A��N𙈌To�N�]�4����;=�P�Л�@�/�(�$v�tj�����a�<zUQ!�� Z������h.��|{阃��k�^��*�������׬i�����dCu��`�(���2U8��=X�/0�����ȱ�!�	�-��"NCk�CXEB��̿��.������������X�p��םׯ��W7g��Gl*4��!BOT���T�2@(
Sobg��C�bb�;9�	}�

k`�X�;ba&�����"mB5?9�x��hЛSi�-�&>�s2�����sn�(�J�O>�l�d�U�J�{dTT�,lY�d�F��v}�Vtr~�hs3}�8�NA�	t�O��z�"]�� &4.�s�2c��Dv�w y���j���r*`&^�v5��|�=�=.�&,����c����O���I���=��22Ӷ�KE��h�,(*�\��x��ʓF���3Kh˲��|Τ�>R7�ĭ ~��~�`ǻ�==6����B�{�`���i{k�D3��F:-��y����[���Bv'�K��9OG�Q�Ԯ�>�j�E$�$��p3�o{�|��-��H^��,���:�ڡ�S��/k�`���H�6w²+�6x�z���\�W��U��w���Ih�5��<[�˔(ό��7�VD���	%C��8�^a�H&�K�#��d���R��6��'3��Ω@�{H�����8	�Qˌ�2�?���XF���(��S������ h�bP�bf�Awz.����ub�ɛQU��� վ�:9;)p�&'��BO �P��qh�Ϫn��8̸�>���&�U����/�� sU*��a�;�]o��}Ub�Tx���-'؇RzF�a���R�^��aσE����k�<6��i��`���O�$�`�M��S�������E���F>�v�Q����I�f�*�n�P�t�������W%T8��á���U��E��m��Ͽ�U\_{l��<_��Q�8�O)�?�7s?}@>o��	vb����-����^Y����������Jr�p�*�xJ������^��_��FX� Z3��R֬{WRS���d�$���G�u�ʶm,P��%�]��8�M<C�������N�ǃ��/)ĭ�e�0aP�UL`��2�d�k�N���9�/�;�Hz����� Ϯ�O4	�xϵY�\�zԈPN�;?�Y�6�L910��uS��x^�ޕ0Yh�(��^��>�`�l��V]�l�:��h7��L�/�uԡf[ҐNCa������@ʹ�l5D�n��6 ͛�}�q=��y0 t�rY�{���׿�À���U.�&dq���E����$RU��5F�*������D��B��^�J��p�iYHS�����1Ơ2Ğ�x��3�l�����^b��gl�#_�G6Y�X[&_0�����x����:�b3Ia.�5�y�	H�*�i�Nپ�~-hI=��۟K�o�JqD�� �8���r]��C�w���#3e<���Ɏ�(�g���ڑ�x}	ر�M$7�����Y@Y��U���T��G�.+����d3�p �yI��&�^ ���M!��C�� ��gU�	6�f�����*%��\� ��ە��r�%M��&��'L�P?�f��7L ��y	.M;Oy,�X
�V�0�-�~�;PS�iM\(he�c{_]�l�p2���,��gܟ���x������:��9���{)��W*K�(���(�f�>�{,9Bu:�y��A�D��3!�?Y�.S���Q������.��T>xa�s:�<|��	�:�n�ϋ(� �,�R?��d:��BH�L[�0�^�/��x�A��0w �"]Ӽy�
�qorslŚC�H��x%�M�K��`U˗�9���PX@�e-��y/8^��0�@Kc�Z����y�J���K3��I�p�u����ԟ�t-��+�{�$�OE��_yJ��`�@~����s��VL.tUw�z���[*פ��P=R�m	6 ~&H\@A�C=U_U_�ϥ�V�F�5�E�DH.?�� %B�Z����'e??h��	�����?���ö<hż�eG�i&�^���5����vv.���A��O9#V���O���s���Wd�.��K��1��(-���аF'��(kD.�~l�Lg=@��7^��?��T9]���bѲ�ĭ!�ޟ/�BG���\fx_�)>�[����Q�Fb�^u���2 �a��A���I��0d�[Q��uo���H�4�3j;Wr\&ǜk$p��U+e�X6�0�!i'���|k,�{V̚����Rm"1"C�T,g0����2gV}����C8�>��(6�m��}�N��@+�!,5X/>���os�_<�� �ws:b`�tp�ݪ�o3b���$���5��[�K��F��JBT����1�k<N���[Mb�a���Wjp{`'f�A�XP]Z��s�h�5G�R��N`Xl2��m�����J�QɒM�"����3]\#�TD����V|7㗾�+��8��f(gK��wY�lզ�j��ټ���Bp��(�
=�d��i���';�zj�K����Ћ������K��b�~�;p��X��k��N��v���d�妹&Z�e��)�����]d�һ�M��6�}T����6I �;��Z'�fw��(��*�22W�S��N^�U�.�{4F�Pr,�2�bːw�v��1�8A��|������'����rR_���:�{73��=0][$��A�X]�=�g�T�#�0U���M�2c����8*4���NP2�<J�o`�`�!�!�]����>�U�$b�q����ӳ*�'Rl9c�UR֯(����Yo�Vجdi�۹ن��|������;'}�ن�����'��<&�H��r�]i��*���� �Jh��`�HW%�<�]>��ط�'����ꄮ���r�6	�.y��PüGC-��P��q�1���i|�k�������|�	�x���S*���!�P+Ń1�hО�Poa1[�� ���Ou~��A۩x�}:{q=ȹ�1����4��s0�N74���U�.�ArvHL����vadt��T�ų�;�U��]|M=�z��
�7XxBsyo�쌪����Q7�+�<����&�wR�Ν��� ��o���Q��=�n�d�0g�@�5Cw�@}��ѽ	Q�M��qiێ�1W��y"gC�N��G�M��s��e�C��[�1@�P��֛�.`�-􌑥�fsF� ������w���5�g�++�jB��V��5�x헧!���px+�3��Ͻ��������7gF��%�H���B�R�|Xwn���4���fm\x���-4{,�t��Q�xhS�ht��	5���$:��ߢ�K�5��ur�,���5P8Yv,����*��J�}x�xS&�R������f/�3K��?��4;�[��H,V&M��ep$����6-���e���}�I��5�!�Jb[�Ir���^�)~b���j$婹�p?�.�˚�^]Pt_��t�����ځH����ȱ��@��b0Ne{�y�n���]���cܓ�E��fH�l�3�p�®h9Z�=���l������2��녔�����dC�4��_��C5wOc����?q�t��	eR&ϙ�:(�ahKu	|K�`��������^�#�����bN��Z7Y���W����-'��N1����|BHـ�+���h�C��|���j��T��_�nR����#ж�r���%�f���|���6�1s�֣�Ɋs���f''Þ\ڛ�D��\!�X��!ۆ�/ʪT	o^��#`�"�|?�8S2/}La��j���d��e֛�7�>$�2���%_۫��m�Ɠ
)�������_��՞@��1@�L�m��o�,僸�4' ?;��>"���43d���yN���6�+����7�s$�7qϤpͩx�)�՚Dhq(�mpSQ���:M*�Z����`�Z$݇JX�{TY\A������B"6� �ߗ��y�1��9S"����*9�W!w��t�G��9��δP�
ʱ���sĜ43J�Ǚ��M�����*z�� �
Ն:ˆD��Nk6�r�#�����́
8,�V�~h$��}DjY1�X���g�a:�K!���OEB\�$ϐP��G>�R$�<V��S�e!�Qu[�=~/�T�۪�ȼ2>��W�m씼�m�])�LKw�������(a��/�o �<ºg�ӑ��ɼ7��1�)��5���<؍����9r��n��︎��D�!Ghk�
���s���J�yNy��?�(����]7n���;�14��Jh���8�MI�� �
�m죢�k@$�³�X���/N؇t8�@By����F��ϊ�ݗ�����O��g+����P�`�����W��{�YC[&Cb��\�d��l��L)U�Mpl�vJ�V���T�b'�����a�ĉW�L*j'Tq����yt�pߨ5�2�ٯ%n>;c�_1'�1S��fk�&W��0|�aiMi�WN	���c������\%����*o��s�ǳ~��cF��ZU�IZż����5iW|}�e'�rm����)��ʁ�@�s���H%�E���[��i7C7&f��a?�&L:���Go,�5��V��]`p��;@['�tc�К��&���L���>2��b|����*aD��)���UN����(��1�=xۅRr��j+�D�G��
��xk�[p�z�|/�g8��~A���[�#H^�����3��+E���ɹTk�7�H��Y9;�hk���o�[̺_���z^�=�I"Q���XJ���U��
������M܉��nɞ/K�~�}��P�֢�&&ZzB��5����$d�U��~_�7\M�Fr[�����z<�Ծ7U�M1�b�cg��	J>xb��Ž���:���D�qW�����n�p�f��}*�W~a��Q��V$��K���R����3�4�0�໫�O�tL�r�Sc�y�x��=+%��ե���K�� v?�όH�.@�"��U����!.-��̧��q��|/P�{xF�"�����_�(��WІ �bq��"0&���<}�r�Y��l�y��Gꤰ�9c��F��n��>=Rk�^����{�q�|\~�]MgO��}���<��mu^tB�Y>Ų��a����P��7��w$��i���@��,O�?.�Բ[D+��%���֙N���<?3�f�J���hI�����Ux��F���'X�c�byx���sHQiN��;Env|u�w���4a��eiŠ]lK��Y�)K�I����/ލ|�q�R��2RR�g�̩���1�z2\~�W�`RR+�UrXR`���M��=����BՁ�~k�����ؐ����N�.t7��$��G4/����q'���ʔ�<��t�wk�n䥶����N6:���m�q>uF,��p���B+&T���8�	Q�|�����o����e�r�B�&W���d�ۙ$:���"T�<qE�%/�T:���c8�:Y�l+j�Vs�e�2ft$��L�eľ�n��-�<�n2
�������?�	}b���JM�o,�95�lE�/y}�$�8�+��b���N���E4�Iu5C�[�H\�c�8�y�!�n��./�"y rs�O:�������@�;/�4N�\;e0���.�kF�q�5N�x����=�a��q������s���qq���i��N�
Y���>}��T[������-�ON�ΠZmr%F�B�B���4W~��zߴQ�I1�2�a��{Ƚa�ݑhwLAjr4}�vd@�̔���yU�7�M�o��%�7���8qM��o���]gW�Ԋ�hBT�Hav�ғ�Ԫ��J�(Yqlf�Q�d��!��1I �=:�HhyT*v��b�r룰�-�SH�>�9&7p�c7�r�m�y����� �w?*!䘢��z�x�@jB�8�H���5k�������&��� Ջ��9�m{��`�!��/Vʸ"��-�$v<29� *��?t������n���`��VT1i��`rAO��g�/U%�4�|��~��`��b�V�0Z�7Q�܂NƐ�/�S:&p��KW�t�.EF�].���V��c�l��E����0\�^�������b&�n��v�C��i�H�*K~#��ܲrˇփo��-�t��	a#��r��O�V�ZNkV��G�[^(K��o/�O)tv�i�����n��_	آl��}"�5�$� �n�'yk蹼&]I3�o��@ ��`�m���������S����^X2�r�K�ǟ��6�8�����#����:���"�����6����iJjRr49�i~8�(�Ĥ�F�&ϼ£ZGV���af���?�ƫ�z=�L�6����Ƨ�>�f��#0��Ϙ���E�E!#�w^������!�֯پU`|yռ�+,k�B��z�Rg-�#۬�iu�Ԙ�xz<h�;�֒j?t�3(>$B��X<5�u�ύ�[.YNq����uL��L)�5��:��pD�3w[�^*�Szv��'^��T��)O|��	�9\
X�EU%����#�����[�ᒪnF�� r:vDѶ~����8�M��a������(�R�GRp�s�r|o����
�6��r��^ONh�#/c��Mn.���l�Xq�e���j֡� ��
i?��3c����Z��\E����s�^,������qB���:�� �D߁)�(4�T��5�R%Ps�f0��vk;�WN�
����p�;ddK�l���}�(�]i�:���.�Hz��W��㗕Jzӳ$'�PbE�C�&ʒ��{�Si��*0���w<�Zqq32-=�6UC�9�̢�r_6�d�
|�9���%�#b;S�i���]aX2 �g�(y�&"���7$
jF(�L��,��u_�.�����ˡ�QhLA��C����)J~E����p�y�G�\natǬ�unw���astc{�'|�I���0��B�������� ���^����:/�%p|���5j����>҅r3���VmS��w|�*76�A��A<ɂ�U�):GxNU�K�?�݅��k:���o�p~�>�!qh�sB�����a�P�� ����ؽ���|���Bg�\�������������OבIѮ� ��cd�e�sn-94*>�t|I	��)�������@U`.�����8#�����h0Z�4�N`��G?(N��;���FZ�¨�t�$�B�ij|�Ϊ˻Z�BOrF��臏�:�T%�����<@}k�#��3��,�&�S!(Mt��� �!��C�.j��ț�m��
!����I&>rѠ�K\����XG���4��Xm|ڌw�y,K�����`dr�J*M�m�C������+R<C;��4yv�zxɅ�B<�/o��r�JM�~=XF �6�Ȳ���v?8��s8
)��U,�>�ޟe��e�y?~"��FyǏ[�-hE�'n����(�LRX:#�8��G���#�Ů7�0�xA=|n��B�"vȢW7a�3���1�ۥ����N��K��,�5��f%�7+&�����+=*���5��͉�B��Y-ͤK�����n����?��).��|9$��[�e���YGp�E���!�T"(���/�_�]���iGO#	�|�и�=wjK���c�u��T_B/`Y5���d��x�4]�L�?]N! }u%"/b8]C��`���`�{���:��Ԕ)�l�_��b�H��rij �-��%m>N�fM������5/����PVG<�yֵ�)��� ���U�k_���v�+�m�J-6�;�͖�i����OD 2���G�f�+��o�o���+肽!���ݹ«�D/M��p9��
T�M]::���S�'���ӈ�[��o� ���s u�&c&���D/�Ӌ��#~��awM8-kA��'�NI���yG�(,�~;F�V3����C�u1}�+{��7���o�w���gj��i,���"ɮ1K�|�z������I��y�B	�����Y�{���}�m��*��`r��3e�Q J��PyUk(�%H�IB=-^�����b���r���$�b��z��o҉��-���D�&-�F���FfY���8�p�E�@���)���1���z˔[�op��ɐ���<�e�?֗-d���> ����Ip��������&]h����+���u�}�5�4�CFݚ�Id�=C�UܓC]_7w�)�SM����Z��`fae)����YB�ǫ� &��_2Ⱦ���w�:2@1�"{���sYPRhɭL�\�5����1�8���v�8��{���čy!� ����bt,��'���A`��D��%,���Eq�1l�9MG���	�7�p@{op�y�����GL����"O�]���@��R(g�x��a�x���P����ā��'�w��Dê�;@�Z�nX��Sպȏ�m�"C�˱RF��C����䘉���U�D�fʲA/ ��W1F�N e��fZ�&Ḑ���]\�թ5ɨ�c-ao��JHF����a�٪��r��UoF�B)�-D-�r��;�/U~Y ����C�Rb?��-��%�. ���*��@g ]���'C񷪃��X��lH��s_��jEń���KތFN"SXS�r[��[���(�Ei;���7iݏ	��ui�Q��6�s&,dP
�|eZ���YP$i܆Q�Y-E	E��F�?�G�f	�[��q�mEŉYI��EC���5��p��VCB��q��n^h��6Eb�Lb�*�Ѷ4��`�J�^�4�5��,���������su�=�}�W��lO�璊TR�`����?��G��b�b���~	h/k|T�q\¾J�b�ѨK��qi��o=��X�m<Ps�۠��� �N|Qr��D��7���¦HT"��[x�v���<;WKٚ
���gf\5�f�K5�.��)$�+:��뒒�����W�P� �6ݧ�}�D��Y���#f�O%�
RU!�q�
HC�7Vi`��V��
���a�®$��@���v���<`�b�ݼ�<�l"|��>:ԅo�r1����r��$-"	���A��[zF�gzhȊ2��*�|B�&Ce+��-�X�7���^�-�y�>���`�:R�"����)�X�@��VW�hMC�C���Grt�,�u��RA��ъ��h������[P�1"��ED�я��4�n��}�Z1�� �t�vzc q�����d}�IHN��*j_0�x��M�AkK�Cs�s'����9F@�î,�e�񟰞τ  [�{ �^�Pi��M�V=�]:�qkOKrBc����ɺ]p]~�Y�w89�x��|D?�.}����_�K�v71L��0��:���/�v��)�M�J5�MD1�<�nv�!Hu@��������Qd��GG��
��;F��A�� �H�o|7�������>���,O�D!���u���?����olU�G��pѶ}�=�κR�O��]�&���>���r���"���9B\΋��W����k�/��ߧ�ȁ���N7�hp��!��tt�����!�Chj����+89�C$��p��[ ���7�Va���cjјMO�������o@i�xђwN��
>������!�5&��|�}jґ�/{L�� 3��{˂L�e�Ӎ�M��Y)��_b�lZw��X��=�fe������N��������DrǥJ2�Eq��p� ���E��b�ܸb������dC�xF秷�O���q�'Eo��et�	5�c� s���V9}���۲ri�v"f��6q�Wqy�"���.a^��������ڏ];�/v,�a����HKl���M p� ��� \�r�r�C���kK�)N�{9ߑ/��ކ���w�d�-)G*	�G���Y�FoH�����/ qO �F&�菼��Øc�u���Lb~��v���,����_R����X|���В��f����/ys�* yg���J=t<<R�"�Ԗ
v�9�R��h�3Z�e+z'[�O�ݘ���E�����y�븣�2%�S�A��=�D��F���iW���V�=��07�N���m�So � �U�����o4k��{`-��*�����G5����I����a�B�G��I	5v>�P�a� ]��G,��m��M� H�k!_���p��˅?�N�M2Ý�SLr�@�Dɮ����DZ
a���C,�`o��ׁ�3c7TA�U����!�nOe|�d�hg
9&,�u����w�	m�sq��}�ܚ%"�}�0��3>d�� 4{�Z�(��d̉�dCR��#<�,/�x�X;�N���&4yi�
�'F��됺�.�I`i�3A�����v�,�l
u@��E�)�G��E�����o&�Լ���̲0�a&9��poV�,�j[���������i��O{����@�w:iB���u�}��zw[�=�P#N���K.َ��Ք�0\dɇ7��R}���s9w�B��a�z-�����q�쉬G'�B.��ZH����'&�Á|�B:�*�?�"IV����?����ܷ����O)f�;�WT�6�݃n<BoFy��Z{��7��O�ub���ɓ�D�
R��ҭ�s`��)���@��!3�"�*�/�4��%:�Մ��0yQ:�E��ڡ���CA���	܅A�b�:gS��
X��X��S��!���L�2�T����5eC����XW^����s|���~�����6��D?�}��q |I�S������kM6��Ҵ��w��'��c(���Y;C�k�R�|�])��ַD�F�	u����Ai����e0v�aR��-h��za��7i��(��;Y{�	��PjҌ.���:q`t��Ԓ�?K���=j���rW�z6C���ۅ���@�����S�:�S��m���B�)F�����e�z�k�@C�b�l9>��]+���x.�O=a��� kG8��,��� Ǭ��r1g�F�'�
�M�T�\K��"�d�/����pz��Lx2��c2�N&O<Oq�*��7Kz�	<�#�@��P�(�.�+�t�òX���ί����밍����5x��Q����k��lZ��RjD>�=J]F�4���h`�c���L��퐼�|����,�cs/�N��[_��?�3�8h�R@Ú�(DS���967_�K<sB"H�}���b~`��#,#4��˙�+����U���]o/+����T��ӻ��C/}�x�|#KC�ug�'0s2j��u���L��n���s�=���=�Of����Za/�/i|�+�$]��{h�G7��*׬.��Cb�h�� #�4��J�D�f$��	�g�nu�t��@�	-��I��R����{pQT�Xȿ���,E��]>r&(j�]��������uA��B>[�4�����ç}).������I��'�;�aojE�jT���� @�T~]V�+��a1� ����,���}VWէ_	?t�[���G�o����l������z+tn���%�L��. D�f1,�~�q���BM��`k���&V&N>*�L7ώ ���|�mz�|~�ufJ�W�$ԋt%�E$p~%J�ˬR�BJ�B �(�R���{�LT�Ǥ��6{ �����H�I!��'5+&]�6!=����&!^��p_�<Z$\�d�����/UҪ��j_c�poj_�z+X�YH)^�X�����o\��9�e�ռVg��U���.�!�d��������3�8��/f|���e�yg'T޺g�<�m�f���`Se>�\�"�R2�,P?b�RՇ/�|7��;-�:0�iI��#1j����2�)UI�^!dx��>?Iς�R�`ۄ|q�o� O��x-)T�'���wd��[{��c˕QZX����ԌZ�K8��~�:��E�T#�E�0 7��i���+����'%�����$t�]	_���)�����D��xu1Z��Lrg~"�d'd`c𜫔�cZW����q(ۇ��Nף�sجAeCm�4Hʜ������[����Ȣ0Gn\���3�K��""�-i��%a�Dj��iր �\Q�Xf�"r�4]���ԍ(�����'>!橘��Cf��qխԊt�-�V�?�˅�:��R1�{����R[�4�`�*>C����wF����jO�ʬԹ/�Z�eO�4Ğ~����_��`���Hmsl���I{�|���a��z�ύ��:�;�K��hv���E�KUj�,i�XpK�����{mb�*�<FR�/��|C�'����;�3���P�c�q��d�N�b�.{J��b�12�޷������c��<A���҆(
|�k��p�Z�:���EN?}��	����5���C��������St�h%vCaz6�
���mtK_����W���kb� ���%�ƞ��^�����߄hIo�pU��ޅ�jH�
�OR�����\���eƣ)"�Q�䧰�M���^�g4�<��ih�f}��j�y6S�^���()�I}u絃���Ow�4��U\�!T��u���dm�)��h_s�F@0u���%6R��D�S¥��3�5�O��]8��WK�t�);�k����{�T�ϖ����[��,��W����^�ַMl[�	8��(o>ɟ8�^q��1j/��mq��m�J�dH����L���]_.hT�>#�ѩ�BO�W��M�^D<8�d��PeS�Q�ǣ�q+���Dc�����
 ci��l�����^����s��cR߻��@�֥ƛIu\�l����x��0��1�|Y�m9 5�������elf6�w%���'��X0�%�PI�R��r�\(��l��N�\���&?�Fa�`�5�З�v�k�|��
��?L��@�h_��o^Z�;)��M��C��"�)�[S��a%���l+�C��J�vB�+�1?Y�^>�ԃA������@��ف~T�a���g:��[��,�o���>v�M�1H���a> M�e@s�mUxw�g5��*Q�j����P�~�K42�5M�ӕ)�����R��Bo����t�p���׬���5gy��|#���V�8����bM�F�R�}�a˔~��"0ȅ�s����1m��r9]��J.{mI����e��ɠt�����Ɍ`�N�m���'6�԰P� &4U8�"+�&�m:�]���?���Q#8����������������-�5AP���tiHYv�-\��yB�~�h�L�Ww�_��yN3QĈJ&?��C�a�O,��Q�fÌpI�D��$�k���z��'��UP�U�}�yv�{Wױu�߷գ��p�s�����ws��yW�ĉ�1�+���#_�/
��S�-O�7Bt���L�n�]�Tv��r48ɶ���9�o7q5�yکv'�n���_BL�
�!JWs�7r�.�#;� �K�Ҳu�΀�����m\U��>�{e���je�Ç��Ύ�Z��~K��2�oe�4��`{���-k$��7x�ciJ�c���^$�p�ԃ1��q�Fǔ)>N�E�0��#�؟��z%�mw�|Ц��2�אq���	�L�eY�t{�/>j��C*OIK��J��nZ^��	.����se������	��q�'�zvw�<��%UH�h�^�%WC7I�|)o>�7V�IR&Q�t��3�*X��`�NX������>g��x:�����%7Ia�M-��Lz=ʆ��� p|�V�S]�?4n�?��Xu�G�����0#Їio�
L/�.H�kp �(%/͞)5�����4�K7YY�/���2�dտE�mR�l�	D`�L$���E�S���%�H���c�F�$5C��V7/cW�&�k�][6	G�����C�6BG�kӷ&P��(�HJ^�+c�4�Rb{�s�����j���f	���R&�7Xw~�v[�x��In�~��j�s�j���/rJ�+�0�<DΛ�eo�&�!�.m$K�IIX�6Ի�,!J\+��f�\␑Y>Z���RǶv��=��0�Ƌ؀�#-�}�2p�S��9��s;�|��Z��4�;n�#����~���� ����s�쪕]��t�q3��p����d$�[A�K���~W��5_�_푇�����.R���̺���7m��=�}�L��с��;?�ժKƃUR�̋Q�s�A7��<��2�g [#�}Z6C`��#!U��`	�Y�x0x���Q�x�H���ծ
ԩ��[��j1e	�Pfp l��<����ɎQ^lA���%d��,df7j>���a���t�N5. ͬ�K$:�S9��� �g��h&ãg�ذR<�5�`�����D&�~f�s��+&Yɞ(�cׁ�鉶Xɓ�h���
>��0���bC	���N7� "��|��
��ǟvp��k_i��I�A�/���#�l�m-�#��q���w�q25��w�P!���z�En�f��&O[(:-���y"�Ϛ�������Ҧ|����_:}wE����ebS��[3NC"�7��뜀}>L����4�^;%����� �{��zF��Y�٦������&YZ<�JO��F���	�%�֥�`B���6�a
f���¿����o^���h��M��f)u�����s��(���?�a����#��ǻ�m�;L���f�̈́V��+.W�Ĵ0�L|��\�a�ݙ�N�ɴ���$�o��}��s3!*�+��i�殬���k�T�S]��8A�W�5�{���u�S�M�r�l�(�Z�6@��_���n .�2��4d�l��\�1pDeJ8�G�24K�&y
[���a2K�B,�|��ipr����m�a���z7 -x�% �u~>�����t/-xc��U	d-��5�����Y�i�jgw��@�[�"|���T��[�<v�X���fd��s1l)K��;9��n���9�����d��7�C���6'k?�M��r>�׵Oh5ˣ��� �}�f}ۮ���e(��}�q~֞�Lܔ�D�ь���*2(�3f)l�E�=�ӷ���r�P��W=٨y��S�(�����Q'`^BA��Y�d6Y[����C�|���4AA�� ��qtM��\f��e�&S�lP�aYb(jM�\X�g�MMT�Hc�t�: �qG#�|��[El�,)W�=qp!�B4*^�����9�f:�ߧol j��^[��v�N�L��L�$V޼ȳ�q�N�u�n�yY�r>$�������l����ƍ� 6���5�ƻ��T-^���U�#��)ז�4���d��	
�����6�����y�\�۩�TUrH����oUG��pށJΘ:��_5!�ϋV�A�/(
���6at�̸�(���J\)��FH��z> }1#j�$l^��ʤ6b�pƩ
��8����S�t��p��6/y~���#s�,�=ԫǗyn��ە�/��Wm\Eh�1����%��2��+Cb(:�凿Dz2�ϒfZ���y����ڪ� j�z�P[o�{4�=�e�ʳ,����[� ����hs���1������s���%��ɐp"�{�����JL[��P��p�(�����$�͋c��@%oBר���ʙ�fn�3�Ѭ0:��*�V��jN��(�j3��gN\�2S���=o�sw��D��W�;g�/�,��d�ep.���gi�2��[���j �N����|�	˲m_�8���lkβ�.��o�������|n��]w�˫~��.7ĩ@���+�'��O�t�q��q�6}���ܤ���Ѫ����9.B�,���������ܘ��������E!D5���ܓ��sf�e�Zl9��RI��!�>W��﬛�&:���'RL9Ij['?1'�lY�rώű]X�d`թ\P�w��u�����
�4~��c��~U��>���>#'�EQ����_".f��W0�21*��x�@w��S}lhp2��$�Y�Hp/��ڼ�@݋��(Z���s�w,�k�<S�� �W\YM�����v5�1���Y#���ܺx�c'ϝ|.�����雮�����+��ì~�y�R��Ƅx��ͥ���i.�²��VV��nt9\��ܠ4�B�p��5�dX`Lt!�'����*Q���E4@[�gw�]:>[�%I�[O��H�� ���8*�c~�t��ԬxI�dd�ع^H����0�[�gXD��_�����gBU_:|e7x���o�����D���6���j!�*
C<�46�az%�d�^�޴ݻ��C�ݻ�`j�9O�v_R&���ќ,��8z�\�Yc<e�6$�9���=�Q�$6;��F۴��=����`�)D��#yʞs%)��o�<���5=�jS�֝y��Q��Q�}�K$�o���P��}bQ�=~,r_s��������h����6v�{���PP�f!�SjWB`FT�?��Z	��7� c\Gb���R�����V2VU��(����D}_	P;�]��L�s���<���fΞ�W�-���S��n�x�.d�@�&=�������X8���)���a�:!��n5�R�<T��"/�+���9������B��O3DP�[��χ�����C%OM�S�ӏa#D˷�W�y��j�\n.{������t�m�^PR�w�/�����y�?o�3���<%y��?n��L���f�4�@W0l�JO}</��A�k�*"��oS|�a�!/ŤS=��tG���..4뇈q��*�#�1�����Hz�GR*Ɇ��a#h�~��K�sS_wЯ?�r��~�nP0�j�B����h-��ss]�����1�:z�v��02��Ӑ�_���V(���)�*���}ƴ��B|B{�}�Ƽ�8Oh{]a1o�`Ժ�sD��|HR.*sP}CB�G�DC�*�R�w���75��l�a1 y|��3�4\��=��tA��;���ko�l�/j�?yG�ܬ�[��gO����є�a�惾�V�V�2��K�X�N��({^m_vo>�W��g�a2��e��F��Vj����Ze1��J�s�G�өIU.�7"V	 ��3�o(������/J�ڧpm>�"�k1�KE���:CSI�en���}y�����h	�P�{SW����!�.RQ�$�;�Yk�Q}�4!������R4�-�æ<�}wU�\�1�^�̌�R�ƪ�vv��~�_s���[�h<E���PR�+KK}[���Ѕ�Ѷe=x�%��#Oy��ɴF�eS]E>�d�d���yVl܌:s6�&��rүN�EHvE��8e�<$��D���w�w=�a[ǯ��䱻�5�U�u�����Mf7��{`&h�n�5�����	�Ys���_�Ld��aȇо�$�E� ��4�j�@�P�&��0V(�����`T�?7��pܤ}[��Q���ڛX.t,�K�B2|��D	IT����	����7<�z����E�=/QS+kwg��
�^�f)93jr����C���+2qMd\�W�Mk�I5e�?�B7L���=
�_R�|uQ����>;�7^����\��<)Q�yHm5��$��?�3t�7������� �h� ����l�P��D�I�05�brοG�T
�ED1ݥ��.Һ+�W>������ �.�zz�KT�r�^��b�1킒���ی��N�`��]�_��9(��\�pa<��(vS[럋2��í��N[��%�G\"yBɎt���k7�����X �n-�{�Ii�g�f8K�޼∰1B��$'�Ge�<j�T�S���-�)>�����7n���ϒZ`R-�g�[
�O07D�F#�d$>�1謤��(�m&x���l�r�'�_��"K{a�=��qgrr�Ɩo�Z+@!��
�^��`�L�4m	�8:�JnFc�L��21�QoJ�W"%�Ӱm{:��wW���T�
B:Ȼ�5������![g`�=R��nB�����Ja3J�Vh��a�2�=���T������*���r��IA�PWJP]��G#͝=!p�WGmw�γo��$����J��'�J9�6�dU��ʂzĎ�_�Y��z�ޜ��	c�_'}�oИ^�/d��]z�P:q�$��{��x� ���ѐ�_��:�hW�nW�=�r���D���e}0v���m��<�\$pُ4dw���]2�Юk"��?-��~�X�_�H�(�qg��bn@t��2~�[W����h�O��=��,V�븉�Ʃ��3z�/�򷛐��0�х���D�?ʴw��@�m��:���#��OG�S�����Γ�fũ�'wz��Z�F��EI��ڕ�e��<�� ���2���}�H�͐��Q��!xi�{�������$��2�_���/��	k&/��0���t�b���ZP���A5��J���x�;0�-�q �"���|��P���Ô����Mx���;��Ҋ�*�(�9ՑB����|�K���U�G�M�����|S�4��Z^��޴R%Gw�T��A �MGW�C��T}� })p�#���ĥ&����K"�J{��W$K��Ą�A�2	�7��1�
.�u��9O6��u���V �Ǳ�^���F.��[���F�C1>�^d!�V�Z��8w��[�6���{�i�ц!o���o�_q��sDb$�F���.���;/���,}ڋO}�O5o��������r{�(>PHJ�	���$�������`/1^֕ڲ��R�L��6�,�q#�뀙�[��q�e_놆������%�	jS�t��;�?�U{�`�8�r�5�:�~�����^��Z &ۇ�=T\�$$��N���V�(��]hsH�u�#�r�Ǚɢe�N1�u�ξ��dA�ݐua�;���@���*��.-�ƾ�p���|�aa#:��7��1�0�	Z2��y�M	����k���Q�p$"��}A�dW���Ǡ�-�ژ��>���+�ke��E0�y����-�U����Ys,'Qp&��vBL^M@��e�W�K�H	�!�t@�F^��YQDT����J=:���z�����[�}�Q�A�v��v:;P$�h�q��:���*d��%s��v����%���x�0ʫ�|Q��Cu����6�j�g�Ƌ���'-���y>�r�łwY]+�q��G^�G��xAi~_������G�|�c��y�@�1;Dh�!�7��ݧ���Z����fH��^3�͕��T5��rd+5��9`}@�^��j�o溺僵��󻠔(lAR��A��i��ڬU�N���YO��C*������|Os���>���&���3�P<�_` ò\��׵'�ڋ�u4�h�ӡ�ʡ�cJH��-�M�~n��w���@��kX|�2s#���|�hm�5_��"����z��ja�����P˪c�G�Jv7�0�쌲<��oF}=Q��kr���Y����tg�"-��{�閦8k��rC-{1h�?��X('G}�. QX�1	�K��<x�=��7c��e��o&38h�(Ƴ�2$���B�6տ�',o�gm�~U�=9g��EI�%���CG� �w4c�l�@�_Q8F2<�F�vI��l�IH� C�\��b�o�_FF1�FZ�Á��a�Aܗ�:W	�L�d��f���+D�3W5�����Z(W�Ϥ; /�uv��UL��e��K���62�� hn���]�(|�_�SNh�!��W!bY�=�x"x�4���+ w��s�"O�'��&I����9U\ cS&�����EMI���� :9*����qE�<�woLl�uc�;K(��<>�3��Z4���d����9��!��J��?��@ե!�����
۞Rx����;�}Qo�d��QdhH��.�`��B1dD��$�<���	�W�!�>EA�:E���t��F)�y���[͈������x˷ �H�j��d�MX�f-��h�#�I�%����v
�FCk��{�_�g#��̩�c4zO��A��^fɃS+W$jm�m�Qtzq��vN����@��T#BQ���h�+��9TxB�Qa��іC*��jY�l�����CQ����������+?a*�y������ ʧ�0M���d��}�|OA��?`��x��aX����oM
vb��ϒ%�d��^o����ٔm҉ʌ��� #$�1_'����D	�|q�h���2"�H�s���́����S�6����Y��۽/�و8H�SQMC[H�B,u���bE�4��|��O:�3Jx�ѕ�|i�Ͱ!/��K�t^�఩BX�U(��퓹���]��9��2,S�6�xU^�C���>9��Q9�4"ɸ�Ɖ2e�)�U���т��g�
R���q�a٥�d��D�\R�y�ۯ������S��6ZfY�`=��1pw�j&��=���g8IV'&U^he����y�*`^����no�N0`UMF��5�c���n5%�Qߔ\��̇s����T	��S�tX\��(�8j�[c>�N���O����vTx�m��D7��]<wPH�#��?�.�I����'��L-�/Կ�Y��dŃ�Ҙ"_�&ZW�'^׈����~�=�Z}v](���V�j��̀ֳ������T 0�C��M���<����"���p���|UxHwd�0vk��y�����{Pt:3�����q8.�������е������.����|X�0
�=�������Z®'\A�q�l��<^Mi4&�B;��Ͼl�$��d0��k_X�Be:��*-���H�s��۳̨�G��q�� 9 E+�P�6�������yGyb����^\��!V*����t�ֵZ�S���eyJ?'����=Ⱥ�=��i'_���]��Z�����HZ���9�~�� �(˔}XC����Eo�S�����E��}L�"I�ۃ#ׁ눿�JsJ�¥��������Mp>� �K�����I�G�:
�eZ�U�s+spmN�Z�rY��%=�F�]#M�W�t����#�	�5$���$k�*b���J����m�]~�iAcCp(F	��bH�q.㷂�N�����һ�I�����/	����OO�!Ղ�Ͼ,.��B��/�	P�S�� ����=��z�<,lS�R?9��;���۰��V%��ު%s����f�Vp��\���'He�4d��6�l�������ӫב�1�X�d��l��F��"+�H85��>�1��b�x�V{�'��&�7����b�T�^Ҋ/$�R8a�҆�ʄ*��T�$��϶�K��H���L#�?�c�zes'?ʑ�^{���?~E�Ǔ�aV0���I���KH���`K��� q�7�
�/Xa�_Tsd�����(��vZ{!���,�D�����1�	[tb�h��P��Y9����)Q�/���Q�~���"d�_�O�*�q1u��e��w��+)0�<�ߥ������/���ja�t=C�r��D����5�} ��^�XTU#�8�1S��Sث�Ba�얋�����-~�77h��Z3�R���Xf=�49���tɹm(u7��J���!�����ձ��k]�a��ߍ3�TJ�#8`wR��v����a$+��T�H���E��l��X1�ӟ/ �5�7wj�Iqy�.S�0'�ث���� C��>��%�/Vq˧�=��xɹ9��Z-�d����!'r~N���V]��d)�y�1i�R>}�ɯ�6�@����
z�WyT�<�7���[���o>�t9f���0�wN(�c`��2�S�&���A�Ћ޳DlW���O�z-u���/�w����Pq���~XKN��?��mؤ	����z�N�������vb9�'<1?Ƽ�TBD����`m�ʴ�L�3d���S��Lo�.)t�e�F�j�L��E	�������"�u�,!���j-�% ������-�s��Yp�o���f)[뿺��vau�^�h��_KJC��u�fLO0;�/�6Z���=���M��KJ�ʞ_|d"5�ܽ���W���=�8�64Q��1N�r���t�^��_O��ex���ƟX���
�H@GM��j.��D=�7�O�����3�x��M�K�}�!��+�#�L��A�Qi�MW�t���	�E^άD�#�`�#���E=e���:��e�S�~NP<8�LU	�P���E5����&��%Ѥ	�8�^��m�X�c�i��g�q��n*���B[)D��f���܉K����D�8.we-.y󐚚�u!���raR�6')8ĳg����%C�0�@30 �Y(U^����ܝ�MF�d�����/�<h�lE�<m}ԟ�_d���
��uE|PM����x�)�ߝa�~��[��eϰ����W�t�gLil+avo�~iQ����~~��������;(�d��YC�艑�h^�$L�0{� ����:-�1\o�!��,�0ηFZ_����F-D��:�-DyTǟUȞ�y'��|�'F=Qh��?=���� �؛�7(�(\���)>����70v���A�t�`��RRQ �Y�y�L�O�� �[j���	����}9��y��W�9T��Cf�<x�����(�iF$��uS����Qp�	by��O�>Ӵx+��4��sÃ�vx���f�ˠ�J�V�)[��cɥ��%A|�] ����AO\�(��=�2l�{=��U�It�3�ۇl�'�JO�tMs���>�v�M}ׇ�!��#�\�f1�ʊ�k���%Z�.~���=5{����V<{���ͻ�j�-$�#t�ޓ�f�Ϳ��8h<$Š��X�����oS�W�!Y�� ��{������}j��H����x�e��`.�a_��]��!���M9d�]�虞`RL�T��VK^\��h7*���5?��&Y�j#�,�X��Nw�����D�~4v���I��(�y)6�so9�����.��` ӣi�v��{�HP��L&!��AW���&�7�>'��[�RY�{�t8�}�B좤�Y�lU�H�H���~c3{~����<ht�\c�s�V ����j��EX��_W]���jWR�'!��K[A�z��}�/�P���]����d�f�v�Q��$8�>�kAK:�?_�u�Tvi��R�Ǳ}`�@/6����m nk ����3����h���O?͖��)7~v�2��a�V�l[����B�-�b%�Pp����#'�A��E[�u?ʖ��(یT�Ҫ�ڬQ����(� Zġ8J���s|U��/��X��dR�D4{W�r��L?�:'Fe��0xT�Xs�y��h�˷@冷�L�[��7[c,J[�g���Q�kZH�Y\���#��q���{Dػo����Uq�J���5��%L�eHܽBIEڀ �M���Ԥ���h��A�c|��8�8L��>^ ���@���������*�_��uO�_�;#���~��8���v�������0\�~�=΂t:a���\�E�+ͬ��v>D���*�F�T�헹W�V:ɏ4�v���JL?m�H@@p׶�xR��q�\�I�(�--��zh�Da0������ڂ�,dZ�f������ i�91��&CUX�>vj�9U&�D�X��{��i %��&�pbrp
�q t+l�\����ۨ��m`X��\��߀/h�ȷ��;�Ձ�fT4��Ĕu���9���!J�$"|���ީѹ]KZ@`�rK�<er��O?�?� d�g>�z�Or��=���r���s��LH\{$1�HNG�s p���=��!b�i��YPe�c�o q�x�w��t��T(�z��h�
"�ȑpub�=�*\��L��!��ճ��D1�m6\^nR��Z�r#�����L��$E�3,y��w��ژ����U|�������/�a����p���Q�f�՚{v[�Fb�L/T��q��u�/������hԩc,��D�}��Wy0":ȕ�i�yM�zG$;�4u�I.%�S��%��wGHk}:�3��������fam^��se
?.�r2֗+E&�K����ȯ���{�c\�W��E��m��P��9�b�B�1�L���M"M"�ji��c<=�|�3ˌ�35q%n �Q�#�d�|�爔�53x5<��Q�#�W Nxx�qM[�#^��6��6|!��H�1PEɂ�փ����]�Q[���]�	egn�)��I������e��	�Qfʤ�q��T	�7<�l��	�yK�3R}a�?E�+�o�%�c���}K�N��s����'�;�Ul�vquV����h!����%�����@�sR兰�K�t�I�́�Fި�t����VO��:jX�"��X��[��o��]�b�{^��kG�e���.I����@�ՠ˂ЬT"�f<=�*f�xq�����i�e.�� �V��N�r�4&J���ͮgTWa����$���2mw���*�F���=��p#pʋ����:+dC6���Z��_2'f
�q+䅥5Q���:7�A�k�ϰ�* ������[�_���z_|�%��^t�����N(��'Z8���.Wݸd"���R
2T�%	�.���٠��4�maſ���ş�}./jp�k�4�Ԇ7�Iv��v?���"�ok�:ɘ������O"�}�ٖ��,�ղq�L�L���s�|Z?��	T_����ӻH�]4���J�Xh�H�O6���Pw/U�>U���v�;R/��B��T�I#��v��eJ�|<(L�.~>=%�cR%c̨w3��!�P]�g��[��I�<-p��a&�{�b�u4�j1*����YCU8�m�ʻ��5Y.C]��r�b)}�K)*�����[1��r���*���� XT|�!	Af-��0�<�g�����c���]�R��%[y�d�zr6^=*QY��S��l�[�=�,�;����LH��b�	�~)�I���AQǲ)x,�T��!�@H+]���:^�ӵf�,ݡo�.b3���,�kU�|����<���,?���0���X�o��Ң�q4�5����(��Q'(��/�Ȇ�aC%��K�UC��:�F�Ux/��ul�m@�"�.���?�e5O�=nz�l����%[�m���R6y@��Q�8*K�S�d:~��O(�����ȶ�ޓ��)*��7�'�v}�o�S'��c|>2!g�
��:�]i��('���P�� 
=�b�1
�)�ڍ���q���ē�q�d��H�К0�����d����Kkƭ'C�Y��D,~cX2�..3�X��8�ݔr�a�7!9<�������E��5xSO�2f�f'�M��F�5�[��P�}݀�6���I|##�4��t&��mO2�n��7�(�bݛ£]��J�����N���U��ن�?���K��:T��S7�&Y�5�	o��w�/�8g[��`���:Y��7�z�o�W�R�.2&��3�\I���l��׸Je�uE��/>�S��t�T��c���)�Z~�� i�:�Jx1GA��r%b{���E�\�FWTI�H��d~�3��B�͖�??I3=��*G�u�T��^���2bU Ġt��^%�I��O���b����m4H��$A��Rc/�f-�#%�V�����H���t0��;�j�;��SBjzG2bQ؋�;Q�ǈۛg*�$�;�ߑ޿�w���⏬B�}��|H�E���&�$d�	�Q.�d��|od׈�¯2��5'�b�8��ؕ;�T��r���Y���Q�"�V��;�^\2��B�Z#=qJT	���hS�\�R��-���v���`+��K9�j���6y��h#�MնIw��=n�7^pFV5Z�/�>dķ���I#�%�V���	��H�,Xd��S@$}a
ʑ\�t�ѣ��|���Q���{D�!�l���̚��A�����,���U�k!3�iͰt�������ps+�*)ˬ���Ö�����3��c�Xv:�`͑4�}����<����l�F9S$��JyO�KuC
�.��f��w"����ʚ�&��	����u��EŜ�4���H�R�դv����_���ԑJ��N���.��bi{�s{yI@�����͇2�
x�b�e�s�?�z��;�B��਒�;��>{��	���h�������('f��ұc��kQ�M�Dk���;XV��a�ͯ���mG�*m���o=����tlA� �f�i�
�u��p��s&u��Y����KR�)�]@��=4X���}�&y��������sD'�t����7V��E=��6A��r��'�̦Թ���S��!p�b�ИE/��ro���e+�O�i=�^��pC8���8�;/ԇ�^M���k��'n�1��"/INc�z��Q����X;��?��Iע]u��Ͽ�Bӡ���Dp
�N�T�����9I������z����ƈ���N>�$�w�6���9%����)����z�����iji�{���V`�z�s	#��v>���b���@�Wg.��hT] ��	3Yɑ��	��P��Z S�t����g��{�N`����90�@��O�3�b/�C��I�u�T�D#G�f�r��?���Xx�������F!��BkD�$�{�jcz��VE���0/yZjcck|xk�- �(��Ԑ�Lo�ѥ#��B�X�>ܞ���_�S�ZV����8�?h��ۍ�Iy�r\k�δ8��z���t7�Q���a����5/����D����mF�3"#���Z� !ܭK+���8|lPTp�2�*dH:�m�`�1p��Ӌ�s��m��nUYc�w����8U2S����S��(I<2S���G,J�u��X������c�s����ϩ�s�hЌ4W�_um��iQ
��埸.g:�^�.{�+-�gZe����S2(il�Bï$-�����N���t�p,(U�;����+��h�)�Z��l�@V���j/�#i�lڃ��$��������57���7y����f�!.z=b͂ ��S�ge>�7��~(]݂��^�bi;_oq���b��m�u�,�*��N��aG���1EK;@y��@8q��yl�uD��� ��b?}��t~���Aum��[�UuEH���P�t�ɶцPu�Cw>:G��%�<��#.s��+�zA�)�˖sLo���v����U��ș����¤j��R�~p�9^U�?	�Z�����
`=���NtN��H�Bfғ�R)vm����8�hG���A5�bK���u�Tol����\���%��*9�����y8�t��Y��_N���T�`��f}�� e�Ñ�m�2�!�D����.G��Aşx�}��Px��eYү�\x5����-5���k�_ַ��<Vg2e��H�T�&������'�\�=̆��j��$�b�\��zyFZ2,`0�j��lUey�>1W9����z�AD習/�����k���}�&(4q,�Ǩ��*�2�O�����O�c *Y���T]YGT��6���@^��� 8ၕ2�,�S@�����w[�C�s/
�����\����8�Z��F_�8�%E��s�Q
�h���:n@ƢL�n+�9�Աy���N��!���6f���:�,�m�П��Ai�c����1�4.K.3[������ZBԇ�7cca&�q�8ɺ��,� 6���.v�o�xպ�)}eQ��26��6R�f�=�#��� �I�su�+Y�	�7�E�Q��4ݝ�
�o����C'��&%�:h�Q���vk\������|�u��>���A�H�8���6S�2����S�`��{�ﺆ�pBW�FҍR~��3y��ə@*��������J�{{�G�:��~���28(���z�S��ɵsқ|��/�9-��	f��!h���mI���O$%$Yj֌��,��^8���<�p��7#5w�N�� �L�ݜ�����_x5�`���7�>�z�W�[xW��֞�%�Q�?GǓޖ���5�cm`�dx��L�7��p�ĸ�Qu
��;'L#w����8"���i2x)F]t���]L�x �6.7A���7�k�odeVmq�� $C��_�	T����]�:���U<�z���%=F@3��{X�OקݣQ<s�
?� b&��
5ۥl@;�5���?�����L�:Bc}S��1���#�Y��v������OY��{˔E�e]���S�'C����iF,�ph�.�� D��+����R������z�F�b�N���:�)�dkA�k�Q��o>�`4N���`x',u�-�G��wҶ��,^K�9�Y�*��p�0����V"
��)���SW�{z�e�I�/��e�;�����nKt�N�şߟ��doTK�� ���<q[�3A��Y�uGVh/��#��pz�AK2��*�l�~�Ep%.�Y�Ӵ�AV�������4�ݶ�L����ʈ�}E�Y���u>{�����&�����`8I��@��F�F�T�Ra����,�ߪ��#���eY���zY�wY�l���'���>��?Xw\A#U���H.e��ڧ�=���²"1�=��ǭ}�JgY�;&�������
�#ѸZ�9��Ď!;��>�!�O9�k�'���і�9?\e��"�xAG��Y�B�m9W|� ^ Hu�v�HbJ��MS�i�s.=O
]��_��S?�1@�AiT!I��'��{��.���o���"e��/��3�w�e�6:q���p�����Ύ�����9RE��&܈���L���5�xH&t3�23�Ay
�X6mXLqվw�S��W1^e/S�h�Cb���_H,�!�,�MKf���S<�m9���A��������>��u�����T��a��^�3���.�#��tUT��ߖ{�=|�L����Ԋ���:�Q郉�kl�8�h��Ȁ��'��]�����C@�|ҏ�6��~5C@�=~����5|{si#�v�˽����%
��]������?;BI����Y���d�r���X 8{h�.ژ�ہ����y�96�݂卵�~^�M�W�K2$ x���w�5E((�_��m����Yz�=��霺[ߩم0��S�r(p �sS"'g
N�%$-�3����9�񖆚m#й���$7j؀]
�E�'��a����rE�=�`*�$��p��>X7`b"���_h�B0��z�B�_~fkPɢ���ꢛ�,�ܛٍ�vB����L�P��5�L�iR�EPg��d0��/��c�FD5RՔqG]��Fk
I:���@�a:t�A3������8=�^o%:a�`�č����w�Yh<���{�&fAi�{�A~*�L�P:{F�ْL��t��]�B�z8]�B��/���Z�y�է���ؘY��ey7B5������jf�$g�'�ov[ 5Y:Te�~��������hcPTd-�6�Ú�X�ځ>�h�v��F�Xu!6�WCU���2ƛ�<��M忸�vB;P�v�O���F������#��/!�y��B츬w�EZa>�k�ؒ¾���.�O/&h���K���QLo��O��\��x�{Ը��4�r��wMoM��+�w��Я쨠k��!:��w�94��x�u ������X<Z$m�Q�bX�H����6�S��X�Vaݛ�툪�
_;�U� �h�X$ ��;�Ҕ�]OF�e�[��z�'��d�@��8"��]6MW������׽b�g�	��L[CC����K&S��������������<�~�DF���OV��q�֞~����`���h��c��^�In���f��jfsI���U��{���G,�XK���=<�>6�XT)$�@�m����Z�"����#��%�7oL����U�ͽ�Phź��� ��ȁ �"���3�����`; Cջ����̲����ٍ/V�>J".R`��.3�3� ���x6��'�؉��]j�T�Op~**έ���0fm�2�U��>sV�H��O�~s�8Qʱڔh_qyZ��~J`��i�W��"�W�7+�����~7��yP�q(]@e�K�t�YKfY��������o�[e�5����r�1���b����v�A栊ԍV�WW��F��k����$����Żc%���xc�j�=���w�����w�yv�aֵ�b���k���6�����H]�A35Wi�N�6lV)�\<}�h _�S���4}���w��'�QD��t�c��z�Gv���o� Qʀ'�nv�j�����Bļ�s�@�b�y�(h�5��7�?�7��ɴtL.����ϱU�&�;�-?J�����<z��D���o�]�����g��'�T��e��M���ǩ,����+�k��*�Dz�:ڢ�x="A��rظ%}������S����h;�L�3�����n0�2���NZ�����b@�*eeSk��į�؛�$�o��<��R�k����P1_�'e�~��ZjW� $ܚz�6���e���vV�λ^%�=���e`��7ح�_�f�RRD8=��W� ��1��j���Pk�N����ÇMK"�4�����l�������vFw��g�����%Ӡs�=W~�����-H9�T��c��iɨz�I|o���+��x�]�����
K�(�M����-��ӽ32�ģ���Q���Ī�a+��q��Tm�ǇB#dY�Q�:C����V���R
��֤�c���b�ŵ�}3!�uњ2�Λ��#�,k=)��K�&�MTM�V0"��5��"Bs����7`3Hux��*�b�X3sp�=~����k�\f~��i& '�����u�d�������XMö�$�*��(�zMrD!��D�]��Nz����� 
>������7��|7��:Y.1����ͱq�V܇w$�ޮ�И�>���m'��O{��� ��P�v�ñ�aE�9r���_�j:�:m����V�\1iݽ_T��q?�:g��k��5lg|,?5��x�*��m�7��v��Y3��|�	���K���� Vp	��J+h�Y朶̗�O��u���˦)Z�y7����Ҧ�W�~�_�����V��0f��J"Vv��f�I�	��Z���,<��cF�ͨ	؁~��G9�E"�����ĕ$T�/�@\��a�j[P�N�ݣ�����:����
M�ԝ�U���h
C�n��x�fEBJ�#�N��N��ԗ?=웰�WV�(j?���8b*���o^F;�t���6)�竓̙'L.������R�Z�,Z�����6Kwȼ�g�H�����Z�����u�����LD���V�(��Q���_�e9R�F���K�����	 �k�0��,��ct��M���d.j��}*�Of���~ި�3{�O���f�!�����9f�a��%�s$cP�?��Z���!9;�q���r0;ֆ˭f=2��Y�X�o�l� ����O4��,_UH�#¢�&�B/�쮂lr��S���	_�l	 |#��I� +S��	�����^-g�0���t�5&��F ��QD����n󥱒���T��.���y��:�E�a6t2��&��=���� /�l�.�n�k�t�7?��a��� B@K^z�m��sy���e��M�ݥ�H���۬���A�)��=$�. `�w^͑�=��(+��ll�؇�Eɮ���}�0�[1jBj��
�y�d
���;�w
zJ�o�a���L'x3%�H��ZtYt.�+V�̂4� !l�i>A�hY����.��ʲH�)�tPָ�_P+ %Ö�����]��X���?pK@p��R�[���O"��hrJ:�?�}厚I�?H>��ژ���	�M�KF]
� �/�3�����Qh��L	���%���=i�Π��k�������I��`�Tqi�����j�x�9; ܚm�0|�� �@�A���*=�藺*H���洶��ԋ,J��'�=����]����'�*�V��č��`��s�	B�X� �.T�R�vJZ����%�so������������fX�Mқ��(>��O���~0��1	~y����:�n���-aέ�yVЦ�g��'�Ì؀=�K���E��������J�B��(t�˃D�^{h��U��{f��>kU�T0na�����(1�/�`���&Ǖ�����9���xo�z=!)��jKCf^�1M;���7��:�=9��Ӌ��5���-�RIކ1�W�w�,'/�4�y�k�p��������(W����_B;��k�DNu�eJ�;[^wj|��)DT�3n���NЊ�y�l�
�2�
*B��
_��gf �(��s�vr��-d�"�׍� �D-K�-+L�֝DU�AV�r�e�}�@q�S���X�"�['Z�Ė��s�1q����M�����$���n5q�n-k���,J~2�i5�"N����=Z\�r��iǈ��t������Ħ%�����:k�й�#�NJ# ����V `����ʱ:F��3G'¹�kߋh�z;���3��5��=-WE�KPB)���d1(��d ��3��t���.08�K��^�q��|�[���F�h���5����
��d��q�߆�V�L1��?�z
7���,��@b���aV�m���*	F�(�����t��t�م�H4����O�B0O�.�Ӿ�״h���,�.?51m�8Q��5��F�Vj��0�{�z,+�9�Iy$S�3�~�vUcޗ �%�0�A�$����{%����O$=�e��ee�0	$��@��T��|�$7��fT3p\��n�*��gB@����/Æ�`��-��`��o��7�x�s�v¢�$62U��Wf��q�ٓ�v$����]�aX1�w��r�WK	�~/C�)[�Q'�Tn���x��>�8 R����Pr��M��4�S� ��S�LѻZ�~i���YSM�9�*�B��>�c�H����
�~�:�,�3���q��Q#a��`I���c���JA���E5*^�ƏiP����G%�7T�덀���_��++�6@)��<�^�|j~g���t�>�B�RF�D�n���{x�� �082�PI��gS�~@v�_X8ᰘ�똸ޥ�e�B���y�⏁M֎8#X饅���I1��ˤw5	���G�@.5���(��{�����KR�]�����C[Un��kN�muR��@=5������c�9&"�^x��'�;����vPu�1ո�7;1��}<eӬ�ť	P���FL������&i��D�"H<�A$X �
�ߞ=�*�w�x��צ�[�wX��X�e��S�f��)Aa��l>F$��	��*
��u[*�'44[L6`�Iҽ<�J;�X�%�L�*�e�^�YCd�Rt�LӰ��!��,M�B̤���7�C��#9���9�̸�?����!�7�n�L��s�)��o��lG�	.��Z��Ͱ7?&v����R��f�y��Z% k���"1Ysa?#K�;XO�ar��E�kC��,��5��5(��9|�7o��Ћ���Ē�����x[�S��m3��̈́�������b}���,���R�Ր(�}�b�"kM|f%�~�[2b��bq��$�Y:{��Y4�1�p��w5��������x �ħ{ѕ�z��zx��r�����1���;
����i~���C%��
�I��4w�E@�GU��ô)g{�kn6���n�V��Jr<pA�	*|#���P�3��Y���P��џҎ(U5�Z9�HZ5�M}>W����q�S>0.�G����dv{v�D���
t��(�kr%N���g�'Vu1m�'�a �����P�Gx��"Q�kC�ư~󁰣 �`3{��@�]wݚO���y\��:sp{~��jt5�@��(����O��ވ��4!qR��%�E����AP�;��Ǒ�7Y�<�6�7�}_9�K�{�����ޟV��^���u}.gߙt�J��W,�Ŧ���ʝ�>6�n�F5�x�����\����C6�+*���$�fb����^(^�F�Q���lS�Dt���-U#�	���i˄� @x�3
J 	��(��3��]z�+s���Җ-�|�A �(��˥d����������B�O�)8ك�披r��۳0��dx��� 4WWI��^~l���:8jG�.�<�Š�BZ�h�C�?���>&��}��piA�m�澐�C7�[ �I����0�O<g�Sw5-@�!��am�=����y�6兪�-�����p�~�	��:�`����K\{R&E�D'�5��D�Ӏ�1c��Pt�k/����09Js�Ǵ*[�`m!=~�${��=j}�P�S�I�p߹ڄ�x0�CB|�ԇU�@G��=�;����k�W:kS����#�)-o���(5��򶄞������jh��*��R�"9$)	f�Х���W�%�!�Ͷ�9L���C�;�,�`*��o>i�����OmA�1��S���;k��>$���s��q�Z�Wz],h�s4�;c�@�L揲�����n������f�ϧ3�S�RS����p�եi
�����H}��]����X�'{'}
��ge��.��Y�lٛT+��y���g[k.T�>�h@�$F(�8S�'�Z��֑u������7��n�����Ԉ��<Ɗ*Ѝ�=&�'��̊k<cѽ�z�D��j3].x0�d�=��|%��J�E�p��lt�~WB�ă(�^#��W�vo��Q�J���	�NN}u.ϼ(�|�V3��������O3�N&̎076�z��'_A��O�ķ��̦H� ^9%��7y���#,�D���ۑK�MNx>Ĵ����D�*�&.�y�-��z��z�8|��w�0~�\�f��SN\�#�C~~����$��^�K�֥��;�l�_��V�m�E�?V�t~٢��Tq���D[\j��NQ�^D4�2[UUKDņ�Ȯي#n���`�Kr���޲q��Ď���q8:�{�V�'�������76���ieK¾&��q��1�:��i$��fɋu.(�P&=���0q�K����x��7Jz�������K��������Ls4� \s��lXB��p�'{�w� �5�T�����@+��=�[꛺\?���8x�����$�LC$�4��C1d�d�� �2-��s�$�Nnn=9��2�lT�#�_��s��#� ��\
�
�w~����@�b!�E0!r����4+o e��(u���p��1'y
BE����T�j��M��X惠 o�F�^�	�.<�w�,� d�+���.^R����&�Zia ����
�Z��@�3��嵕
��@z����i�������yGU���^�쀹��lc���qZ�&G�k;�,�C�D_f8.�]�y+@�/�>��9o%S�������+Ƀ����絽؋���]�,7���S��J'\��;��aK"���i,5���.��u��0/#3k厤��,�^��wݻS��={�1q�,d��,Vi�mL2�&U�^�{�-(ou�.���d�Z2ݟc���sĶ��~#\��f�M��yK��;������50i�A4��^��G�V@oi�iD���wD�@�'W�D݁/<읉m&j�H�[�#R�<#x�m��� aT�j�����)��-Ѯ�c���޿����ph���>�"�*��#���md �	���A������w !�	�=�hٓ,滦7>G���>�DCfhaJ�|H�y�V��F�,`Xf$e���[0Q�ۣ�=�V�g-�;8�^��뫌�>��Tln���ˍ����Fj}�R�`���w'[��3?:d3D\O��k�N��?U���˗;qn���fL������Ox�}�^��B�d�p�+�͋���jG�XLf��AYX�[��b�����;QC�Q�-��2V
�0+9�z+o�p:?���7T�:�����g��5E^
��B)�/�(��u�t7b��AE]=�߷ߔ{Տ��-�<Q1��~I)��f^)}�͔��wV)�}�^j�GV͘�Y�a�%C�(#�˛���u+j��
�ƙ���g��k�kC�H��> �_ek�� ����^�"�� hε��^eʲ��f��N�d2�h���."�^���q��� ٓ�Y��~�Kzp3T��M��S�m�8��[\.�!�s�&"�����:I'ށ_a�����ˀ�Ϸ<Z�-w�ৰW!o{�=�Z	��Y�1�`jbղ���4�N}#�/��c�<��)���Ks{��F�L��p����0�P���<��h���f:=� �ձûy�`aJ��Yi�'�L��X�SR���е�IE�*Չ�j�	I�7�D��U��ӽ��U��_��!94$/�`I���L�uR�����#җy	�|�u	�A}h'G�~.|�g2ı篲cv� ��G���;�w�Nx+HM�����gō�Zioh�3�ŕӃ���.F�:�#�cr�����1���$��O�q���ΕO�WY��w�Ƕ��d
$&��(#k){�F�QH�]�c��П�6�ew�˄;<*�Y3Lg���ޏ���{ÿ�'���
�.⿽�g�S;�_(�5{W��4n`�mS3�]�Q8��b��:?��	�
�͹�;�WݞUa<Q�2b�_�+����M�w��䩌������n� ����=�(;1��h�暽Åd���澢tj����F����	|��P�h*��[Z��"<��H�dPr��o.���F	��d��k�n����]{�x��Y��A�*���R4��\�W��.��UM7��`6���vXO����2fd!���j����i���S��8�y:)��(~pK���"|x}81�D�^/�dgT�r�c��]I���Kp<m�)|�Q�Y �ޘރ��o�I}�҄5�ˇ��m^��{Z�,�
+���Y%W��smm�MoQ����%�>�r��vP��O9S2C�!F����]뚫5�^�S�d��b�d�y5�1sٶ��C���rƏ��2Vj2��K@�M�W���_RJ��tZ�+=#���Ew��VD@��0���\V�/���Pw u��-z����������dkT�PF��!���"4x�C���	�NT����X� 0&�Y�B߽�F�P�
!�h7�̷sW3-KQ4dH���I��f
�U��s��@����2|��0k����i�?}<� ]���bN6�v��.'��=L���u^����4���/N���=�_�'XTU�!F����冪=q;��L�� �V;�̧�|��nC�'�1%:1��W��A5�����Qi�ٱ�B�zF�%*d&����d�nX�Z�b���Bӊ��pPQ��`����X�=����{&>r�6����#^��֯� Rq�Ԕ�j��Ų��Uf���H�fۮ�!7������q|0AX��o�B�U$C:������˹A�H�� #v�]�Y8檪�x֭dM�P�~��.��zb^MQ%�w6������]���<60�^�歙'"�҇Χo�to���&�4�>�U�~���iV��v`��1Z�>E�:���S~X������^D��?�rL�x�6�qCp.�{E!����=�K��?�+�&Q��WZ��*�*�,s��@��D<ۘ	�kC�+^�࿎�<�ψ���WKY�<T���߻	5q���3���A\��ֳ�E�JSQ�1o��߶7�Q�9���o����
���G��x:8g�v�7IqZ|�q�R���Z��ЋD'9�(�����VA�0R\$�P��/pB�*���d���n��j����#�����$���4�د"��u��A����(RT����ݛ��ݕw��`��+�2X�Y�E�*����OdWo���GޛP�gMWB��ؗ�|��¬c!^yOJez�k�#(��^����w*���y����P�	�ෳ�����I��	%d�sx�f.�B�_lIb�*�doJ�w���G�`�}�'G �:p�wgrp>"Ӂ?�R��_6R/ŤW%�A�wҚǫO��'���=��.�K�R���2Q�>��V�N�9ƾQ��]q��W�����;���Y���
��(��B���xS��꺌|=I� $7a;��A�n�N�<Y�O�Fr�T�i8��~����%��Gh�$�RNrĮ �\Ã)O�KCo5��,ӈ�ecT9�D\&���H(�c��ȁ��.]Ӳ�An�dC ���@�/�c����v����@��X� �l���49Lz �[AxO��@F_,� �b?�� �CThN���[����6�T�Ux ����G!,��=|=�D���|%�ԁ��wdEx�=^�a�Bck�>.jB�@�>���C"�>���t�PCG{4����m"�M�����ھ��vB}^�������Gȩ�}Rs!v ˲���C���Q=R�4��]��P�Q�Z&��j�����z��D�ԘƠ����j��Y(��Ԣ���xϔS7d�q2�U��oLC����}f[ze��ۛ���aĊ�m�����`(��}^̡��P��_��+u�}Z�#ф�3���u�(�{�>qH�<��~bU�<Ɩ�4��=��_�"/)k*u2�H�[�ἕ-���ҫ�"0�Nq)֔�?֔T��yNִ#�_�ѦBܑ�f��d�X,%�� ,��	E!��P��_�X�(B�����m��}��'�-wY!w4�����Ih���u��~��m-�%�x=+~���Q��3^@ij���|Ul�%��M�2"�N�8���2鞕�4�E�:�q)�alm�z¯OC��]����ǎ�o�����Dy{�<9�xK2-�
�r'���<�Y|��9^��c�����7�3
A(����U�8��LK�L�q_m��0�#\�f
��!�ƚn�F�3��_a|[�I�*FZ-��C�W,�7���=� �qgD��	.>J���_!�A��d1�j\�����U�yE�6�f=��j��!�7/�����	^t�95@u��_�3�ݕ1�]���ұ&W�����%�M����+���K�Đ/ܼ=�M��#TM���]RL
9I��y��vh���M�.U.�F��,�@���clp�|`����W����N+��/���+�v�k�4�cO��6p�	����(e2{\�蜳��l)pE��*������B4쟁�홉<����4�
PLE&��F���2��m��d4��M�ό{et3̭�	>�+)fR��g�a�D'<7�Ǎ G�����`�I��4JT�� k�n�{��r�m�z�߳nnufKr��?1e%G��:��n��h�U|�����0m��!R���)\��k���P�M/[
�'�ʙ�ᮝӵ���W�[���;�g�I{H���_����%b*tÍJ�@��Ο:�����47��bP�9��қDX]jh@�2�����c�>>ں{�4`�C²	��E�&�ɢN6@<kD���S^�{�!e�V�>-�,DƁ�_���"#�m �?�!)�עC�<q����������d�AT�|�.�%�(����Ժ�=ν�D���`w�8"�����@���޼m�����Cck����WG<O|P'&\�FCwaBʅ�qz���~�F��І�~*R���C����D�u��ǣ�Y� �O>Rz��>�L/C���jw�Ǜ}A��)�m��X��Y��9�%3e�w
t�5�'|^A���eL*� �>\I�R(s��N�X8��N�7����q| fa�oW�����
�J\��,脽���/V{O��$�o�Y�&��(�L�n�W�~�Y�b6�'��$��a�ڣӕb[��j�B�V�D�_*���Fh]��6m��O)5�د%�~���[�	�Ϗ#݆�ݶ�(F���h�:���D+�]:ZR�[6�޹�)������WvO��  m�,8�4o���c>�5p�ˡU$É@|�sA�������G��:<�29�\�~�eĬP
��ԓ�{���U�m��@��2,�gJ�J=H{(~Bds��z���; ����իr��"����ʐ]���.P�S����k$�$����м�,
��{��+�=���E/�=V��X0�2յ�7M?�'^n}��c��d�m�&i�-E�|	0\o6�Y�� ���8-�/�zh'7���&	__����T����v�2fB~k+��5`�����z�}f��&ZjU����{�*��w��5v^�
4��sQw��*�-X�_�0-�U����G�~'"�y��C�$�Y`~1����/�����*�	�������!7�6���G�����Ǉ�ײ��¥5���
������Xy�p��є��:q�n'���9���� �:b�?���C�7�Z�b0��ᮒxt�n���}�Crʦ~{�H�1
�p�O�w��U�Ȳ�O�bH4��+ur�����X����b�X�y]Z�b=��/�HݣL����8�9+I�\&�3�����qR�z\�bҙ���v�x���+'iL�P��tÔ��8`5�h~0��yBq��D_�L���́��i�>z	�Mw�:���(�R�M��H�1���xwk�2.G5g�Ihn��Xcn,8|�Re�a�m۟��H7܊��~�����Z�!�Z�4~��툁Ht�/��O�J�2>�4O_���=��u�3��T�5j�A\�w�|�?��^ܧ�Ρ��"��F�|�⬼�/�{K���WO;+�1�3��7��)giS���1J3�˅.�R�(j�Vg/.9���wəj�}���k��< ��S]�2�����>j�eA��N��cw�ySN�KKR�@�4��g��dJ�6�l[i�>�eQ3S'�m$휙��C/g�����s��-�=Q����,�I�X�إD���2�s�P�� �;�".0��h@�}E� q',,�H�no���S�ᶕ�;�0�0]�y�
h&ZX�C�t(�^� #�->�9�h�%s�*��- �o�����U����6T*I��悡��%��KyJ�h���9F�����l�k" ��[ٺfLov�
0yjf@a£���j�%fs�T���b��T��镧
Ց��ubo2������y�%��H:�غ���皶��K�E6v\=Յ��h��Me���s���W���s~�F�{,��f�%��&�E��T����D(�Y�x�4�l�$��F#��@���tw������+��<��@"d��l�����S�ʈ)����'�i�����l�,t��Ȥ�Ù�L�%`C�J���j-_�� ]Q\.i*+���A��+|���)��?�����Q��k�u���q�b������	�
#m�ec�
YBpS��G{4��B.�F|'�t�^�Ai�$�un�`B��q���7�(�S�AN(���![O&d���#�D6p�X^Q�{o�z��\���3�e�"Jr`�Z��,h��:����AR�oa5���2��\0����B��6�=7Ɋ�Ut��{v�>uQ݋N��Ba�{��4����^7�������3�a�6 ��N�%_���v���cG��Y�4c>k�1�s:�.`�D�Ж�Y*�9%Ƃ+��0%�s]⸦$��P�9\/��Ž2$��<l	����烦�`�c���n�u#<v3�_�U�� ��@�m}	:������p�#�"-&˕��z�:���댉$]��k�S����׳���β���A�(�Qx�l�2ۈ�/c�D�75�^,���o�NG�z�K��U�B���>N'@m�����3*�����s?.5��w���w���e�,���.�%/Zҩ�'��$�t�o_�;�K����y�Q�D~���K�@u9]�z7�;����v���Z+/�ޡ�3�^��z��q�kXY���&�r���Y}�a9�i�4�sX��\Rǐl�����p���e�!�͔��t��(��Hf�������y�0�h|`;I����Dl��+��0j�)3R̩�!�#������Y�%�TA��;جEn�7�Z!-:�q�4�}�x��D*L���Qzvj~O��֏�E�5ж���ʠɈG^��@���N\<Z���JH�vU���STg&�(.Q�[rC���-'��.����ŷ�B�Pܼ�ۀ�%o��ҿE���h1������ˇT����@)�,��z4x���eaWM�z3��Ι�Z�Ƌ��:Ci�����Ls0��~����r�]q8���c�qY��F�k����Uԭ�l��ᴫ`%���J��y��V ��&��xY����F]�E�yI�jlכ�W`t����7���U��I2������&/��c���8�	;�bM?�����2f~r��`+����XI��R<�3R	>ߊ��������`�:���B]s�bc���&TF�<�-�6�a8�+=m8�m���=@�Tk�Ce�h���OW��}��h�h�|uL�����2�!�Z�����W��ͱ!;o�U���[@$�TK!K�YpE��9ԉ�L���HK��6N��E�H��Y1�t���	V�^�[{��_���u���R�yi��^�Zy�Mƨ�7<�|�sR���ۿ���w�K.����C,�ר����G4������7�&h��E �|��pYf�K$�s}DQs�Ha=�G�9H'�p������ l��-��r-���z�^���;,#Y�,���4�8�H]�T�fK�����d�s�o9$��f��13�'�V\�-����y1�-gZ��ɋ3`����~����e��0����[����dS��^9ޟ��g�w&t0\B�'/��r��Ǽc�x�ԛ?�Uvz�� ��dLLQ�AQ;ї��O��UȪ��C{ֈ�Y�i=���M�FyQjؼ�����Í,5��ìО�_��P�+�@c@3��B
�0?�'�e$͈|[�}fA�Ųu���u5ܴO/f�h���j�.�M 4�:��t���� 7�ǹ߶�!ƽ�Z6���-B�U��`�-?��z�[��En�^�o�HI�`v��!%�d���
�	��W)D����%�W�3/16;P��������4�N����<�W��8��!�-!��%��1���'�{��|HWd�X�@~R�z��j�s�D�&]p��H�U~��M+Y ���{��Nv%�m�,���^��b�B� ���}#���S�$������$���-#�&S�,*/9��w헕�b�mEea�������	p�J/h�^�� ����&"�ۨ��N��o�?.����k���F���h��r�h��!Pw�2��mB^�'��]�����h^�C'r&�8b��$��?P��t�M�$�����hSF�:�X�S��B��|[GΎg���|M�	/k?���P7�4~Φ��(_J~�l�1.��*�9����T��v9�����z��蘬�č�x@m�Y-aɶJ��H2���Lp��x4Ȫ���8�O�c��z��vhv�z�2fK4����Լ�C=�d�N�7ҧ�Q1	2��y��hU*\��ʐL1�D��*n�5��il� ;H��p@����Ez2�J$�*	LSI���LJ�י]��eM���I�J}�P��i�����?2��س f�a4�.	��n/��ϯ��硃B�D�,ݯ����]YX��Spk���)�[n�^�S�7ڥ��J��[Al��Z0�,�hN[���`�괜-�2�`K��S	)؃�5�s ���<�o�Hl��oM�wd��}�-�У�g�}���(�����
��������b.39>���hl|BȒ�L�:q���y�;v]
%�w[|`�D�ռO�U��^3ns3.�;)�iY����B1j
�d�_:g5���V�b�K��3?��������4�]m�)�7b:����d�#X6�Ò���Vب=o7�@��F����f�^��8�j%��Mvs�1&���ui�_���uK+j1�G�ݓTe����I�!Qn�������R��� ��x����@��Q�y�;��r8
��-���,��_"X
Od�E�*J��H��"9��_���y�t�a�UH��q=~u��8>�hċ� ^҃mb�@l��YW~�!�o�g����(\`�Q�uv��s��ӆ�V��h0��Y툝��`�Z(�`���,�4��[�y�{�-��B�<]��2�}�4r�թ�/�ۧ�m��H�e;�a3[��(9��[��-��y�o�;	1��?��D` � F����A��OyN��z���.B� z�IP�*u�X���:|�ṹ0�����n'��Q�`C�f;C�b��Ь���̌T[���ع9vgS L1�8Wׂ<���
�"��9Z>���o�$A/q,�-kH\�O����pZ�X����w~�[����y����l�v6-�?X9�q�{w�L���1�'
��v�|�,l,���cY�Ƨ5�=K��/a���d/:)�e�imY��a(���M+a�E�g��߷�N+�>[ﰃ(g2�KR���(u��q�X�R	�R�\��7��UmZ����[A�(��(�G��?yBN���0�jD.	�������?��]�3�ޛ�}b��<�(���BG;�P1��r��|�i���j�H4Ľ}�Zi����������|-��:��/�W�Ԃ?��\'+&62Q��}�2��F�V�s��s �N��sF-b����5O�v��C��GD�A���	����
���p�@G�a"�؎��]?Icg��}�!x&�W*��Y#۞[9�9�2�*�-�/-q�E�@W� 1V����l/��
��ӱt��Z2��Y�#����z�j�Z߽e�B��!��A��rA�N���⃏n�%�>�s&"k�+���<��BN���!�Pfݩ9h&��s�E�x�mr#I�ՙ��� {�׊�x�%,�Ja�E!h0(�$��E<a[�?I��Q�r�$���'���Yj��;8�� i`BbRC�A�=�ytQ�{�y���D��B�6�n�O��z�Z\{��K�����ws\{>|#29|�ו/{�Y��+s����L��	�Um����y�Ë2�wyc[wt�7D�>iL�q�RS�<7Md�1����}-$��}*C�XI?ʜY���A����J�t?5�拋��,��+��
ZeD�d`H
�Ε+u���ط���f`��S��S{E��<V-����䓾ہlԟ���06K7	����vH 
�;�Ԩ��w�:�s�t-LE�(O��]'=� �V��}G\�/�P�U �~����F�{�79�U�����n�w[����B�{e$��%�f�L���Xї!�{�,�+�"wDr5���
����>���Nl4������������A��^B���(?�P�Ⱥ�9���zX�p�Y�Cf_0���_��X�U�%���	t���VE��8^TwC�4��z��`��<��K}���a�,-���H�Vta,yQ\�桝*K"S�z]���d^
�ڞ�K�#��J�j�N�N��O����U�T��kv�q���g;���W�y!�ԓ]�7՞���rY�820	QG�(�泞J�����0KRvjQ�[7eD�H��F������<�j��a��`p���k��(7x�W%i�Mfe�x�3BH��_���5��b%�HG�������T'[D�F*$�D�$�(U�P�i�����)��w'y~ܚ մ��<GJ�f��(E�����p%ա�@�\�"F� \lI�>�ڷ�����9���=�ǘJ��_��۹�0�>���Y�����q���`��O�/���U+�W%�J����V���3�7�;c94��Jrt��aK����4bՏ���l����2t�as�?_6W�5��?\n���|��	��oY2��K����6TI~�����!����W	L�1 �yB�&�|�Q,��ɣ�xdߒ���1���.[���f>�G	��������~-�وR�q2�1wQ�gxxc�&m�����9d����Pt'�q��j�:3��]e�x���?���,wF4t)ٲ:�*�]��L��M����#2���~B&�X2�W��-$��D�P�)@��Ġv�m�|��vgF�G�fr�f5E�+�<P���,d]P��d�D���K�U������]S�ӑ���,�}����L�`ݳ�+�=f�2�v�����$������!�N����d|��x���'Dg������Q�ʋ	�i�|�c�l�9�Y���0pϦ���ƨ���5k��c95"�xU�tVsM����	H��NPu�.��C����'�u�-K ��!SL�m�_��8�'<�~s:S�]��^�c�mL,O��G��g��r�_%<׊[��ܧ���*�=D���k����Cl~��݀�%�����5i�Q��� �ݭơ%��N ���@���ӿ�n�tȄH��㤯��]���4�[43�Y��Dǽ�+;'2�g[zv��`w(��J��|��w�!�q���v��t!/�e���I@��ي��#��>:���p���nb-vg\Z��"��H����.[���E�'~D��V�+?S���ʽ� ��6QQ(��vI�eA���/���e�L�
��1� �b�VφK�ƙ�t5�Ί(����A���V�ㅍOO�e�:��YDE@���7G�����;Zw�;(�Ba%\���F6�K�� UG��m1���\�ʦ+lO���Ot�fއ��?gr#�"R��膇��e��K��s�����fऒ��|Di�Pc6az�>��4:~u��0Vb�t��$�&hMͣr�.@�&�}�`�����0S4��!
 �����݃��xk�*�e�-����|ۀ�Utؽ�+�h�DH�e�{�)Y=����	��Z�T��L�A4Ô��:�3�,�J���V�;��_��Ve;yU��	�EFPlX����g��u�����w@����{��6�TH�&�H����9Y�
���_<j=�l�kL�<r&L��Z;꡵��%?:*bmX��%}������i�[;�V�iQ4BSw"MShpvVyK	���r+�N�����p�sc�ԋ��l�l�[������(4.��r���ٹ����&���$;᫮�L-�b�-:�""M�Z_��;�Rlg����A�G-�u����F�Ն�a���;��qWGE��K�y�I�UQJ_���Ҵ�u՛��1q�!�yM�ӥ���Q�ym}k4�:^Ͱ�8':�Έ�m���[�H����kj��{�OdJ������89o��{�U�q��G�~	�:Ӡ���� p��󇡃zyY�N]T�ƛ\0�,Ym�e�?X{ä�{�����b�S��y�y:�
9�Y�wcR;���RY����>e�Xzۂ��"�fP��<�R`���K�F�����v���վ�	%�ŷ"�z����UR�ԉ�|ء$�X��8�3�W�>|�D5��e���-B�U�����q�j��� Jf���z%��!tQ�)�lQ��:uܘM��N��,�jAO�t�T����M�\U7�� v����P斌�E&����{J�$�1��֏�F�Sx��)�S�C�[(�ve/N(����k`"Y~�25d�3�����ct��Lh��ZY��#�	���������Y�c�܀���>O1��2��S�	�rS��d�H$,J�t/���E+�-3�"�յ͊��~�G����+5]�v��s�V�v��
+��Ⴟ@c#�\�����|�
�o��_�dQ���MO�� �B�ˡ�ǈ�A�','%E���@���%��>���$Hb�}*����X�;>F?��.�>�z6�CI���Q̥��F���g�s��0qo���%���\֒hO���5�K(���f��O.����k�G!g�?�L�,j��g������jeQ
�Ϧ���?��
����^�w���$+�����y^읃$�*������p�Rp)�k_$�r��	Ԉ$&��
b�{&ϔ�M{���1�ZSP�"��l�$p�O� ��sÑA'��L���Y�:ದ��Q��P�;-a�]j�<;��XP}�^(�ܠL�����b��]��]� 0�����wǴ;��Ȉ��H{�Ε�f����a=7�8����E�:��:o�p�p'�`X/������L1+�4��cy���	��[ma@ɉ�J�+v�s`�~)�H���G��ɓ�!}��#��+�za90�:i��fk��B�|��î���r��T=/�x��ǿ�vҴ1�����\�!�G��2�F��<ɰd�i�k��1�6������;�\��mj4�v�����:���T�u����� ���-Α�Q���%(oB�j�"z�U���'/ˌd�ϞX4���D�bI�<<,G[/Q����ɾ���̞�6xTL	��f��kU�%˞~�������9��7�*� ������@�'Ӵ32'	�Waib�ɻk^FrAN��X�?�/y��I��?t�TM`�xw�O�X&�T֖�R��.�XT�^;���<nu����@��;�S�-�.�����Au��)�)"Z=��^��R#ԇU{y��,q�BL��1�z�%|�},Th��I�
S;ٻ��H�����K)�V�W�q��j�6�H��(Kŭ��a9�rOܝ�/�uW>H �sm�E��|,�5N����ʼW�g
�G���b`=��x�ָWr�Z����,���HI�F,@��b�tʨ�N4x6�P������r�� 	�,s�={?k�OŌ�>,�p <c�vx�rU������:��^VYaֺ@�l�/@�����%7:��{�.w�q��z��?����`~x]��񋣮C�57_UL�g���Mv�N~i��LGŗ֖���_=V�C��2	����m�����H������m����~:��Om�Exv�'�����H��)��~R�ջB��EV�+��-ŝK�l�55�^�Ed]a�,�`[��hR"tJ2�Q�� @w�e����l	�^x;�(?lַ��`󖋵ګR}�� �ZL��pO�.�;����K��D�a1��%��Nm`\:pf��O��)����J�#YpF��l�'��%Y�@j���j(���:H�T΀��T0�Q�o��G�꾄/ӳ�_��	�����cDsz��Gau�ê���Z-fO�\�]FK����\�Ƹ�M���(صU��*��I�R����k]`;zUZ��r�Gu�h�7�0�}D4��E(�~�e" �rK'���)�ڌ^3d&-4��CbH.���'����@���O7`���3�8�V���&�;1Q&��I�i���������h�������0݋�5,J�O��:�&��YaP���s\��b�P3%H�t-_{},�9��@���j��б۸g�|Z��a��\6�)�ğ��u��xI��a��yy5�] �T�N�E�b_<��1x��c�>��fx$�6�p�/7p:)xRY�Ku�+xN�Ep���C���T!�e7P�������@�əP�z�m@�aZ��!����s g�J�e<c�_�:���Ɤ�S�e���5X��Mi���8�T��v��Q���L��p���:������i����H����'����V�h�2��x&�&���K
H8��\K�%E^.��t��*QzQ<@RCuh�Mu'uy��{ @�;Ձ�T
D�σ�_���㼵O�jU��*��ݻ��-��;C�!e5��w�4�P�Y��<x�곦�b9U�mk!�׉�D	��l�6p�\�Z6>�G=�-���x�eG�O�MyGi�*�G����!E��̐k�N���L�����>�*�Ä}�� �T����o���0j��V�.�[��6��/�����r	i{V�E�e���%�h���q:BK�D��4wf�&ƼT����}l��`~�`��t����r�)_��5Uۚ�e8��`�$��\6�hԖF�gYՕ~���䆑4��j>��pǹ40���z���[��Χ�ӅBm?��H>�y�F��f���Fq���~�Oq�B�P���窮�W��gaP�G�c�ϥ��wo�cP۪G��q|�r���ᦸ	|�u�B�(�?�d��;q���@U4���^��4M�����w�V�ilB��F����$�i�I���x�"$�(��9 ��dњv<��RJ�Ї|�)+���:5ǤLp�N�M�P_��q3���~�?~H��O���jc�����i�.�,��&S�n=�G:dbnV�5��e����d\}��Kb��G��M������oX@�F8��<[H�(H(�ZXOl�JDE�{7����8D@��H@��CؠWqgΙ`�`��=���DL��k����]B{N�q�`�G����]�{�����y�.��Ҏ��+��%��Wa��p�#���A��W@�ʱ��Zy�A�{�F}�]__Z�����bj\G��_����
Ʌ�Z��Muq�B��7��1v3U�V�JBWQw�V�|�]s�~}KFT�<�76�����I}I�H�|;(�YCE�ÅjfH��H)l,�6
<����0�Zb���1�(#��X>��㩹a�R��7;��_�<��pǚ
��Z���)$��5m̢���UN���YKy{��n��f�j	j�E���F&j�0ܼ^��+T��zvg�r�KEz��İ�q��	|fx�hI�m��Na��@'GE]�%�Dk΅{L@��2��5az��A�Yg&g��A��5�Ī�?J���7�qԅ&�C`ز a𷫺[�_ΩK�`����d�7�b
oa�$:�])Js컲�m
���p��*L/dT�k��&��N����1�2;�0U�"�`8�@��a�̐�!�+hL�Y}S�ed���-f&��9Q��B\y�n��.���4Rlx��@�ݰ�\�Ɣz��h�%V�m�C���T�������ݜ��^Ԛ��γVMeVxV5p��I<���
���^���Ry;C�j
�u�V�ǵ)�G�rz<:�{� �Z8Я�8L`Ċ̜�i���{��tA�7�VM�M/+$���DW�����k��jY�if�oDP���dB��ȍWN��&9���H�͞(�.�3Ӥ��Z���o_V}��a�f�ap�ư�ϙ<�#JUq�h����2zqi� uK�5��J1�_�JzZ��l.�3m�OB���x /�R�&��o�_��NNM���]4�g@�f�\'��DeD�19��|p2'ր��q��T�E(96k��S}�v�mG,F��Qυ�<%�"�ҵp��6�0`�����x�zfj�U/����I�Fe���q����#���e��`��)��I�E�Oz���@:��ǀmC��'�X&�i�OP��R�"�6�B>m�;�~l�t�W��I��A��&��!��)��{w�#�l�� �(�����h� D3����+��Qj�����IN�YL�.@/��*���e��̻
�{*;��o5��0q�<뎡t���h=�%�Hh���>��l/�t�l���#��߶
L�'���H��&��'t����Ka��WH�[oj����=A��j��>�o�[1 �x�I�F����;#����L�?5Oߴ�p�V<2*gJ;�j<�л]��<�f p┥���������Q�m�;H�R~p]KQ�H��'nت1��b�|��JDzI2%�X��ک�w�g1:Y�FZΌӄH�a-r���T��q7V�uX�b�Xx�Y_S�������H��>s�$�x���s�Q8�����=YW��x�I��Sc|*;T4����f���{c;��s
��>��L2鉚��-"t�G�����Q�&�A�{�̮�y#n3�����7_����%�����P@��=�;�n��D��&m�?t[Sn�����E���4cU�O��\f-�\ �ZN�?�=;VM�S}��y��$&�� 5�Ims�p���O|,8��*(V��=.:��$W=i2���P�A���0��f�c�O�+�ϙ#�k�!A!3�]���uuAK�7�Vz{tG�SPB��}9\��1?=�+����g���2/gs�$�C����E4��*��:�$�'L����	�Rã�6������ىF�B:s/�2b2���w�eϳ��ͯ��N�%���"F���2����/��d�F�^}(g�u�u8IJ�\״�BH��A�&��pQ�<B�9xܓj�tSg�ٚ%/!�����D+���oR3����r�Z!��$�h��قRPzQ�j��ݙ3�Zw��N�ג^m��yo��0�<�A���g��;����q��&�ױ}Ǖ�S&����j��R1�C0& ����x ~9E�9
7�^}f�<���~�{�Q#��^V�ʆډ�p��tf�%^�d�=?��?�������A�3����!٩XU5�퍝?���ҿ�I�o�� ���*����9(����f�^lP?���[�F,'��UޡcUE��x�P����K�GnZ.҆�bY�V�o؎>��[^Ftt�4��ة<�Rx��,��D��_.��1&˲	�Jo��{��$�tCu��Xn���?q����Uq=��'�$g��2��5jy�#B6��IH��,���M���ఝW�Z�Aس�Y�����	��u�q@�����ube��J��a�:/����gx�M�@�g�ow�-S��6�$���=����[��Z~g���Q�wH�S=�_�'��+�A�����z��s.�>v�t���3�R���U�/*�/�ҥ�ji�:�rû���>����o�N������@Ϯ2�j�wS.�^�	���>/߉�j̿�<�G���H�+U�EO7�s9�����AP�0"�E%b6X�3����-�������\��|f�*\�n&T�F��b� ,�K��K+D��<x�A�+���_���3�[�2�I4���]�iz�`1g�����.�t6����V0�t�-͒�� MUq¨�v��/��|^㌺@�0�y�$�>$�O������{���8o_F@���������UD�;������!��E�;��C�n-`AP�����v����̒%34�i�R]h�Z�&<����}��0$���̡�s��.�lfQa�jlރ��_�Ow�r����g�K#��дV�%��RR��z�y6�z�*#�鴼]U����.�n�|Ep侓��/
\��+��<V��pZ},H鯁����/c�
�37��_D*aq��/Ir�v��r�'[�h��/F֖���8����|�#�M��T�ʨ�l�U�F�qOH�ť�첀�W-#��]����,9�6���R��ʃ ���Mé��-���&��B�g�=�6c�Yu��ߌ����U�@���fIZe[�E�X��Ky��Dfkaz�a��  �h(�����ނ��%l�2Y�IY�:=|�e`�s�ny.A�(�lZHu
�?�X�&��[-�]�j����6���.:��?~����t1�
�э__�z���>�>����4Rf��L��r��g>�jP������4�ǂi
z�r��Uw��i�����-�_k}(ZG<'���Q|���#v$�[��8[˚%�T���Z7��mk:�*H�8�MR����"N�s݅�=ϟ3>Yj��'��&�
J�>z<T��w�^�h�7Nͭ=k�����e����![K���2��$���Ʋ���*�A���9<�[m��-KN��hT������]��@S��A�g]XJ=b�lQ�p'�@�>0�p8g&�{��$�p�VOA�6�Ȁ0MP�zc�z6�g@�[LQ�(+T���c��1جhC�O�TBh��vS�q���z�\��l��u��;���+,�܎^���������rk_E�0�*��5���ӕ�?�]����~yn���;$4�1�E�g�'m�,��~�	rD4
 ;9����k�HRb>#��)I<�c����z:�ĩL�X�(��y���Q��4�ܣ�(�pa6ú�N�uJ�@`��zr��� D�
�'<IS�;(r�M�a%�CŦ����6���ԆЙ�z��[2ȡa�����JS
�i)�������!1ff�ax|�PV_p:4m�$T��m`��yP`\����Z�P{��{�ȯn��g��/�o���,be��op?ϭ:�q�5Y߃�o5C�z�]E�ʩ�����-}�>�	٩�Z����Zao	�έ�0�� Ť�=�ߏ$Q��n�ȋ1��d��r�T5�r�`�YH@o��i$qjF��̥8���/m�d���tl�Z��X6����녇�ˏd��a[o��phg��Ӯ�C��[pv���m���/L��7��{��m̨&U$6b�3nlE�a�+�[�|���o1j㲂um��(#]	P��H�f�f�b���a��^���IQFN�����{D�T�E�d�>��	c�'��A��#���M5�O�o�3C��X�b���Z�^*��5_#�ԙ��ͧ��ae���Ci�����EJ���-U�$���߮�=��#t�h"W�J�t(+�i.0���	ݗf���W8�HTMՆ�ʅk� 3k��@]%������ک��:/ʶe��%�d��e�6�u�El�>C6�"��_��T��$�e����5����Uj���d~�uL�<\�͗��P0���ݢ�U��R���GD��Q��'Aje!�� ��q��v�tÀ�z�<ޘ�DI��U�37<���i�~��� (l�C
]tƵ��Q�Cu�l�t6����Y�`�1w;!�6�6��� ��[�O�6?q�u���^f�Kv����p(��_����7i���1��=t��^�s�`�q�Q�wW��G,��͋3,�N���㦉2qJ�&Ҥ�ܵ�[��ǫn����o|��/V�!�&�C�Pu1����߫C$T��|�i��X��R�+u��%���x��9�yٗ	����b��՟w�;�d�Q{������]yZ�S�Nꙸ)҉�r�9	��P'�\��|����1�S��c!3��e�cƏ����A ��Eކ��g2������m��__���R� ��n�`@����hU2v�CRj8$�\����%;��/��%��D�����>U���b��KY�C ����k�Z��a�&�@�ʃp%ʑ۬>e��}��S���R"LQ�?�.�/�H~'�X<g�����ۛ������i ,�T��6_����oZh挷��~��(i%�@Ra`r[R�T�sK[� �W�d;=Μ�^��8tÊ>��EZ	t��,<{����@�H��<`�E����Y2�퓷&��J g
OC��]�}sSwx��~'ͨ����ф��!�`��C/��d��QL,��3��b�di���S\�֮�ٮ�)��J-��8�GS�d�����Lcf����F�5��+@�u�Q/�-̋r�p���]* �b���@v�_@�����x�p<-dE�j_���i�\U%4=�.�Xe|��*�yn�b�"�Ÿ��=��.�Y_�P�ћA���Ge�t��1����v\�HqzeB���sl"N��dz��v�_���+^���\5��1H�$�=���z[3Q�#,���M�Ơ�:<�^��=�y���\X� �en����o�
:��(����-�_L<��vC�D��./���kґ��kb�ԯ��l]C�H�P��a�|�}N�13g�~���Uz�շf̔]��G��DȔ\+\ �X��c^N�y��V{����	KԯA�|}���*��Xs�n߫l;��f��3��忠�M�}�W�on@wHE�[���C�߻�R�����Z���_�y��C�#��zi���x��bg�RBeє׫�y�	u����'׬��͞v:��i~.� �&(L]|��&Zs��';�d��$��
��oE�)���::�IQ8S��#�GX�t?.�?KFl��x?Zi�1v�k��u�o��,��o2��O7��D��lȜ��%����YFw�b���v�2Ҹ9���-�uv���eR%IA�!�]cc!8���5�,s�b�'��������GVƵ�[���10�I�z]��q��'d�!e�Y�<VR�Ǖu�ܲ�Q���c�-�g�Ħ"�|�0��^�q�B��c�2�>�'�T�9"�w*�T��44�/	��U�`��Þ��|r��6/}�|~�w�J��o�ۭ3O����
��fvi�O���"d&0"��	@),ݐ.o\�����t���=�M>`W��F����8��h�š�!]�.hM�_0������6�������\��Ė��Y�M�l���FQ2��)"��z�M�OL�jv�b�`�O���ݚ,�ލt쓊��Nb
����Ȇb_��Ŋ��uB���^e{�TX��$�E���)<�-{~[�N�VR/�1ؽ�.��R]h{2����Z��3C���s��C����);Rz�R�W�d����68N���W5z�k��w� ݝ;���Kgr�B���s�b{tȫwDh&>���\�-��'��P�<���@���m o2R��\���jo��M�Ўr7�NĚ����4�6�O��~�Ly$1��5��'ǣ8/ ��l���%�h�`��-�1&�txEQ��3#�#��呧ō��{@;S� �"K�qj�@d�V�8���)���xz��!	��N1���h~ѽ����h��E~��`�L�=��5#ٕ�l�.A�ȭ�V-V�=��RT�[EO{B���HHQ�̊�gV���i�@iQ���}`�N��pV4���k���]� �mO�3Z?ʳ���"?Qs&��Z�@ԃ=���7�lЃ�C�T>�� P����`q����Ѻ�/�4��4�2���ϙ� ����*���6��7��*;C&㲁WX^Xb",vF͔%.�����c��Û;�ѵI���(卢�O�M���;X��~|3���ȸ��F�D9��whL���9AG&����5_C��1o��˯3S?F�oA31|%�14w�<u�~�8�M�
�A�+\�B�B�%c+���$	+`���y��D8���Q�.�oI�~G�\����7ۘ3sؤ$gm;й�v����$�e4D��eP��+*��~^�q��b�{2'���]8���Ҝ�ѡ{Y�����ǢM������
ԩ;2��0��?L�r8
�!����,g�w�A��GF廳�AI9����\�H�a;G0/I��m�7<�K���v�J&(�T�o��.��~�#�n�o��%Y�l�i��ȡgvZOpe���)Ks�1-����6��'v"��L�'W�/ĥ���:�%�(��Ԋ�����W�tB��aΧT1Ql�x��d�?��s�y8Ē:�T�)VO�����O���=���p��@A?�#�ʣ�V����݋�-s��u�{�s�X{8�:{�:'�*Vf�檠-73�����|�D�!G4qs�2(!i�R���D���t���aR�<�k�LQ{%ī�:�����S����{|�V�!;�.����󬏯��u�hT`<Z�F�� ɴ	~��NC�$<��d=AW��0���"�Ēd+
pQ_ `
kVu������/�%)X��uI�b.q�6�\'(��:�l�q1K�CA^J��e�I��R�i:�6�Z��U����������2&^���})��\+Z�ˈ���b-(�~k#�Q�9W3�Ai�쯍c/R�B�޵�"�ava!BQ�w���"�єpZu�AXmt�ЖFF7�qaͪ�R�#0�^���[�J<���F��z��P!�K�G��a�S+���u�PE�.�v��cbh�,,���G"ڎ�l��V���$S�KWn�����*���>L�^et]ց��h���a*p��M�Tw���m�b�Un1��$��.�1���>�@"�nS ��G�X�Uǈ�*?�4�3|w�D�WV��?��P���z���5�o.џ��xl忑���y�	�)�n�
�J������
O���TV��]��K;&��`$S8	��/�X9��Y�}���^P��.�E�8r�5'��F-j�>�<	�}3�&$o�(J����'Bx])S���?���N�9����|>������gE%a��q4���mRVi��$S(�d�[�/������-��jS�N,�j��kѐhڲ�8w��:�r �,h��!'9/b�]������/l�����!l|ү�[��W1$��|*�~�;��ҷ"�E�2���M�GFCn�4)�ƿ3�����eYLW��O��t�.+`Ŗ�<��1O�`�wr� �_���S:��*e�X@�h�R)��w��t1�n aEaA2��`�W��D.Nn䪠<,�U��)%��%�z7Ni��a�W�]�J���p���[/��`¹�qx�N���ΐn^�	�US�o1��d�^��O>G��֊��)w�I�'/�	�me�����7Mj��|��6���Ј��s�d�*s��]�0F���e�ܑ�B3*m+л�W�}�#��('�k=Z��f<h��?ml�(�t�0�d1D\kZ �X��<���a�Ȼ�F�璦9��nM3]~m7\K�Rr����W��q^�;�x�v8�����2˓��yi���]X�1�����Nj�C�|�_�/��ɻdk���d��~���\�a��5��o� �W�˃�;��ej�V	l��R��
�U��Zc�K�����9���+�'�W����x��9u���*�1��T6|����R:+�6���г��Ǽ�F�/gE8鏳}C�; ���m`FcYp�aĳ�t�m�<��Dk��]�@5�;��Y��8)4=���5��w	��d���'�,��ĉ�����I
RH�#7rm3{9����n�pRꕢ����͈eކJ�0�J���.�j�=υ�w���u�#rf���]�b�!���� Ȑ��i1J�s��ڣJ���H���ՙ� �*,a����D�[����q_9`�J^*�v��񞢮q��%���v���4H%w9�� =��E�4U���Gf�Jw���҆=X�XZ���,0���R��:��^����@�_$��c}<n��ȶ�s�g8�R����ho��YGGB?��x��83Y	�v�a5�,l�=ۓ��0���q��kOU��4�.1���8���N2���>�̱x�v/~�z,l	���	��F�o]WOw�����r���9��˘2�p�2Fh��M2��D#�ʻ!�x�E���� �/=�Ӵ�����;��Tf1P7O��z��概�y�}��e;�t~+Y�+�}���kl�_
0�	��ͤB��58pW���~�K�b	�+� X7bI�����Y��Q����b�֕���~���4<$)K��D�	��v�����b� ���?����G��5F9���MV�]e��1y��i�M�����\M��^uF-5�H6g�z��_"�[�(��B�<'��q�5��o��"j�kFS�䷫��?��[���c��致���[���ֹ)�܆|$�	E���Zw���5�0��F�k���h�Z��%��1�k���F(��r�çm�i�fm�������j'	� 	�3�~9T5BW���ȿ�ϣ9¶	MN{�Օ��d�+[)!��|+��Ţ5�i��k����/�`,�&���DY�(��L�y��������f��g���q��Y���-(g�}z�47Ǹ���;y�P�
�n�SAL^�BQ���9�4�����cd��6��mo�(eA��D4�����4�^����!�;!�N(^HĮ���%���	ż�at*�q�P�82����"���fMkxV�)�?~x�����a¡�&�o8ca�E9�|��@3rz�ʤ]��7�Q,��;��>��G�챋v�}�8�@@�1:���%<4ĸڦ���j:|R����c�2S%&E;�I5y�U�v�Ӡ�K�aW�� �\�%��Pn�6��c�����GU�jr$p.p�A�ai��C��<Q�H��W���t���[턋	"��?R��j����=�SM�%-�0���u���nS&�鎛�P9G�?�j��1!:��b9���f7����>��@�����Խ�9��2UU5�a@viu��b(CRO�g�<�[d�]� �E+�yu�@,L�x��.J��F��Ó�&[�'_t�-�Jdze9�*�܈�i�G#,�U^AY�V�^
����e��K���Ge�Ţ-��A��jg�u�M�8?/(�%��E���P�����E$|����� Z��5e���}�m�1��E��)��iD����9��x�БF���bp_*��_&d���\�1�9�,��Ȑ1��4����R���be����H0e�艨f��j��9mK���nZD�e+��҄ՙ�@�{~RFBm�_6�}-���G6U�<��xe�\����k��g\眢-�7 �gb�T��/���������U�sY�s$2O|:���~X\v��d�!�I��U��&�%�P���l�P9�6Z�k����2��K���)V���x磕@kS��>zɸ��t(�(���ܭ$ժ�AO�?[W���%Ep����P���ා$EO��&�r��?��a��Û�R?%���<�{���[�6ӱ���:�D�?L� �MqXh+B�����_�+�E��	?��M=��Cv���|��ć���4@�-�_�4�?�����1��w5\Ҳg�E��h��u;3�����O�V(N˼��T�j�Es���K�Q���b=z���^=�><h~m���l���*��~� Y����D��cZ�kr0���SnCu���B���쏿����ǰ{��PvA,I)Yp�oD��~f���W� ���<@��Q���i?�9!��t>l
;��ĉ�u���Ю��0�|����U++�CRDj����ek�E{�EI/�Tm@2IR{���u$�T��l>��4#��"�5詠g+r��Ń�$TeS�"�m�)��s��� x�f�tP�
k$��i.���Ҥ��\#�`��飷��W?���|#d�H�B!�0dk0�L�U/��lA3���1�\&{?ٰ���\�����:�Sn�U~t�)���='�eQ���,�Yc_]�3���%�5~:��q��&a�i-u E(�xź��R&��l������R�10Xf�������MJ��d��oy����5���L<��D���9�ٙ	eO�e:e�ӂ��H��Ae�$©�"���G�g�������U_DBU��2J0qX�9�):;�=(Uj�L�f��C2�H�,�|fπ�f�i�~�9Mz��~W���@�tJ���qok+5^�C�<�tZ����4�d~O]���N�u�����u�Ma+�]F�U�\_.<z~���lR����@w��~�w��%պ`�$�왨ԜNGp�Ā������l;ة��3c6�ՒNj�`��Mh8��|�Ԥ�2������G��,�#	��_%w�!���3���)���F��j���!���I�*x^ܱ�����b���8�LD�C�����l����ɑ^�T�m
l�]�O���u��穾�h�`�R ������(��z��y+��մ���w�O._�`E�(/�G3�^��b���CQ�A�r�~�&H欜��%S>We��d�lV����H��jٗ6�ߚD�˹��t�]a���V���"*��G�3�!��7�U���,��T��݊p>���?��Z���Q֧mt�s+%.���C��\���X���0�v>3�|`�UE���SJq��F�g\�	��A67�{.�"�|�� ��҈	���T�.�R|�j�W��`�z�z&ҧJH���T�'2:� ¶[L|�޳sk/]���c�֋�DV+��Z`�Ў�.�7,� �|f���oZD�WU��'S
S�X��[j�Meu�ܟk? ��͉R[:kG�A��wlA\>V��oߺ���-$��u�LH�쩖q�8�?������L
�Ņ����?������#� �X�A4&#�[��O��w�b�S�c�zy@'�Bn���0�)t�f�� ���s����w�Fꛤ"��dKR�T:�&�����Ql!�ةZ�'=kZ,�����t�����9tƮ�^���TEfL�͍$�&%S�?$��݃�s(��z�ï�:��5zp��9��[�5u���y��W\RCӍ�j��qp&XA"]-��] S6��j�Uԓ�`�Snj8XP��x+.)%�����ʱ��H&>e�
����^W��ݸ�H��R�*=Y��폘���?��xg�9���M�<I��]��Ȝ����J���RA�6=�P��S�5�V�>y]��/�8���u����qmWY�Ģ`�/"$SO;�wn��W�t��V�rz�d6�z��4v]���	��+�=0(sR�w�X��(~$Vs������៕~:�@���y�s,��P�i��PH��d�b�9Ju�� �J�IuT�	Мu̗Ճ����g��.���~T����h�Wn72�]�2���'wE9�@�7�GgE� �s�i�{+:��uVۍ�R���0���ʜn%�|LƏ���lι����C�Zi\5�_��N�w6E5��K�j��R�@�Қ}u�a>���Z��H;���#mD �k;N~4sW�]ġ��S�y7�͝�Ő�(�%dZ�,#tg1@V��6��}�@\(u��VVP��t���o��}8o���R��[P��q�=Fv��7/�_�~M��R������g"��h.�E��q���_��Y����Q^\h=3h^f�P4=�ͱ�9!pg�E> Xq�W@ZB4ě���$$��1�O^C'ņMBaS>j����.�����s'�&�4����@	W�uV�{K���V|�s��0꧌@p�M�}��A�Ž��+_��*��J��>)���/!���Ȼ����$���H{L!�]:��\Ɨe��7����Pg���T.��_.%?�ʯxbu��?5����m�,
aph�����4�����(��7��hg��ޭnh�;!O����l���}yr��@	p�3_�T���p���<���s rG�e���@�Qq1��&��'��6�k�?��(��]�f�/ ׾]�YH�J�q�~�_���^�aϙM�'1�+Ӳ�3!�|C��-����l�3
eF��G�s���|T,��_u�QW7Iݯ�Eo!��.7c��� �Iɼ뫩���~���3H�*�f�Pk�= ���]]^4KI���&**ɞ��C�����|^"�����3C0yX�VF�)�|(�S��6g�G�G�Ɩ��E$@�ӷ�G=�F��ؔ����E�n[a� d��ct���fcf�z��2P
��a���dhz��Ey��a�3�X���0r E,W!��byG����A�˻[VleA�a���!"�����h�N�hȚ���{�NmF~����=)-B]�W���a��f3��+��n`�l�5m�QĨ$�4�^�!����2�NG�>�*���Ƙ�0X{A:��3/��������G?1�7]��b���='6�$���{1�)M9�~$�="��&��S:�%�s���hG�?����3�6b�������1�#�8��ؚXЄ/L(_-�c���fb�B.��NӸ�e�(�E[�6(��f3���F����F��_I�(����%����Ň̉����}p.�NE�L�p��5?��V������ �1H��+�:.���Z��L'�������f����9���O��+�ב�e8��f��x^/ʿ|�j���3$��WOq@�/�v{`���NA>e�r|<���#8��'.�Rq:R ��tR��]���"@�_�h���v9aN�8�F|�1����ϓ��,��B߂������o6!�G��QT�,��灦�p�?V{(�Ŝ_�m3(v�m���i��=ɻ��˖�R�Q�;K ��xb�,&:�bPb��l�d)G*�܄�[G�yZ: zD�	{Bò���voJ,�<�^щcMG���Y4�ax_O�1Iݿ�z�l9�c�$cW`j�nU�!��y5�q��мW9�/~�*J��*��+��I&�;�L�RV��$�/%�n���d~�N����Poi}�����7_8��~��87"t���PUu�ڤbɊI�}ݕܾ�yg�Ȝ�:e��2#�����|�O �+�b}��Y��Ja[����������ml�_�L��O뜬�-nE��Sm�~����;�0q@fD����(�od�(��Y�.��$5?�Z2�_�e���mS%Q9#&j�9{�y�"h�}()ؤ&X�dŠ qi��G��f{��)��Z>�����jF�a�'f��t�hG�YR�w�5ˏ�u@L����w�����FUL��/�χ���H���0��<$�T�
䎁"R+/p-�����(w���LN�?���F�}^7���^o'��,�+
H]���gQ������t���M�d��ӯ����rrE;R ��w��j�
�f��o�L����Ĥ[R���xT)�w�Ƒ�p�N�yo�Eih&	k�~��괅}�v�RN����2߀::�Z2����k�A�,�EDK���n@��6�dp���x]IEs"V��a��3�S�N��e�7�1�MĴy���>gӬ�@Q�Z^H����r|�!�&Bl���X?j��M���ԭ��U�{GV��C~�����t���l�.�z��gV���`��J��Z�L \�Qe"b��CL��m:r����G�)�7��jT�r꥝�T������H��S��d��#�֐5$�z���:���$흫��1c�S'O%_���F^�+TB���)y��w	Pe7����mJ����)ꋲ��P��P�1���J��T�F�d�]: 6:��H|�f��&��(\�T2��I�<Ƣw���� &6|j�K㻗-H�
��'x$8*mM�n^\�uoz��X�:�P��=��"� �]�}��Z`ġ��YI��>f�����d+�vQ���v�H�U�ʹ�~��]X"���8�H���Q�V2��T��{K�K�>h�2�!� ��7�U h�d'k�l����CQ�H��X#���V0�2Ճh��!�b�q����$,�uhwn魲l�,Ń���)΍�"��U��}n���h��ըC�xW�&z��:fǔ)��Y�h=��֮���AD��X�
_�'�1��x|7�z$�,�XM#���t,z�3qVqR�Z�CdM�0�fx�
gqT�e}��lr�p3ӣ�_GL�3���w2U���%�&�p7�|�����o����|�����A0Et�+��J4R}B�r[#��E���:p���}ś.P�Z�����Bh 9Ĩ9}JzTZW5�E��[)7�.�
 ����9SF,��2���-�,�ˀ
+g1F8�b���b�s�^��(:��W��]��c2Tj@g�{N$^*<!��Pv�J�Dn4�9x��@�tA|GH�>�Zs�m�K�4�f�y����dS�sv��J�-�<�/��'�JyN�nOj�C�,ɞ��I�*�zѲ,6I_���&�[�j��/0��<%ٕ�V�5z�W�:�=Td�Qݴ�J����s���n܂�`V�|&��B,�B�VS"8#�4��F�g�҉�ܪ�6v���:�?���X'h���zS
��� �[���� �����'�/	��4xcܨ�Mg���K��74��{��[F��Ve�L�Nun�h4���3Ee3��H$�D��2�G�#	����:?���[�i#����Su]��a��2��@
���4�3S���x��.�|��TBغ��̎;�\Aߺ�QĨf�w\Xm���5b������.D�ң/uC�٨V��	!�@z?�RW���&��X1|�����D��N�Wt��R�Yxbл��d[�[�Mv��b�I<��;�ǎ\�)�Ͳ�VL��/�50+�%sv#<��Q��JY���Q�=
�|��d��	��=I}#����Y���d|I�`+2��T��t���zO}����^�O*1�ǔQ��?,¯"��:������g�8Ǿ�&�f��D�� ]���T����z8����[CR�*Q��Fa�R�O�Kk�J~$e�
n��^ �޳�ԑ��L��!; 	�Y%q&��)�Fs �~����s�!~��\�����lmݍ����#섎.�g��J�Iܛ@AO�)�-Cg����SE�'���j ��1��e4jf��y����]Tg�b������֏�3���Ԛ�-�&���LF:dWNAĢ����e����1	K��B&�⤏�=ڧ���8��o��s��^��a��8Nx}ט�$'d;odZVu�F��k�������a������w�Q���j�@�=.g��b����C��߹6��T!�$	[q����L�an.��*�;Fً�Ƶ�9��{�,k'�3[pRs�ɚY"v�Hb���7��/� ���3{���cf&�-�:���Sl�6���F��V��QK�?��=�^�%�M*���c��v��;hBb2*�7�Ek�Yb&/��H�����@��/���P��-���vH@��ţ���_��O�秛���sN�]� �(�[n��X����w����a�+�sYz���  ���8�eF�q�����
����̨Q�a����=�����۝BU{�����:9�E���i~!��[.��'�8���lY#Y P��@�Yc�,����Q�h��*�(	������-pu��_�9gFq�lK=*��2{�摀zC-aR'�PZ?��U�Z.W��]{S9�t��3!A8�#[㴝A*\T��{^�΁J��%B:Ƌ�b&[�䷙�9�Û��N6 ׭�a|�V�$Opa�`z��K
n�Y����|��H"�)V�0'V��R|���h�5�k�O c���d4/6n
1(�o�>t��TM�i�s/�T^ 5�q�[cJ��P(�0���ʫ|��FW�7��ֶN\p�l&U�PU��aщ������0i"2v�#�!cFQ�t�Y���h�#���Qb4�E%�g]rH��,8 S.1����n�J�.M�<�H���M+߁4��}	s�����Zjk�M-��S�_��|r�o�W�@�	�y�w�-��P�g���cג�vf����h����Q��5��j�I듑^�J�&�*�7�>�v�T�������ۈ�=���|5���Xk ��%��x}֕�*a��[���f���W�x-��'K��qG޸-�V5���-�-��r��Y|2f���ƨ�>m
��r,G�ϻFX����f��J���Q�hl�.1"���r�NFq�Y�rݳ�L\m.Ě��0Ih�Ma�ȳ���:��l�U�UU����
��̠�Q�Y�C����Eׇe뮙O�zrJX��!"���|%�k���ڱ���i/�;�@�5���3g�B�e�u	7������~���XdLJ�✲ү�T�Z�L������	�c�^�q�Jd�H>�z�>q͍�˭f�:f"k�z�������x�$`�0�y�3�� :f|I�6��2O��j�׏��;�����x}4�a�o���gq'>�\i��m���B�d(IثW��ޣ�"������.�̲�q,�۳�\;�KE��hK�l�Xp��'�N�v/�hDk���^%a�5�Y������גq����x0K��&i;��{���9N�n�1T����`��ʻ0Ks1]�6U6���V�K�����H~p'��m�1���i������j�)��͗ן�q1��ʏ��R_�ΰ1�=�/�n�&$p�,:�����YtmSQ�}�@<�*����-�����x���W�9<�|��6�_�LK ��m�!A5xC5����"��	=�F�!��Zj�U\�3��|�}���>4�U�>=�>S�uA��:�Fg�����!
+��43��ɖn��<�>I�uF��.�10�����"2|�ۛ�I��Hx�t�� 񆤻��)�'�9,u��ʉ3�\�����I|I�̉.��s&��c�	���n�X"�Ů�QSW�`h?`�U:w:��z��,�C{|OJ(S_�!����]�v	̖��;$]��oW�fAn��{֏s�������h47K5tj���a�B�c`�L9��|.�_��D>��<%��3�>ND]Gr�0�1��^��VO��
�֕1�5��ĤA�lh�ڎ��]����̝4]������8cM���G����`ܡ�`�&�J-SP� �	�p8y>� =��J�=˔S��7�D)�(��ң�JNua����wo$�PS��
s���|J���D��Z#w]l�9zu�L���Đ輥���FD���ѯ�n0���zJz�
)���yYU4OV��7�S�\�	{����}��i˹a�������-w#�X��A��X�8�l��%�0�w����CL	3v�Q�$��������l:�d�R�ؿ�h��=�뻇O� ��p0F��'��~��@�+!
��K��l�J-ZJ�S�?�/i{�ь�G|�j�F��`�ɽ��"�"����Y���)�^�-���s&@�IF�]�2{\a\q�ϣ�ý�65Pj��`z�h+=�d�H�g	j��d������U�m��]�>'v�F�Xu�Н��EѬĆ�ƥ�>�Q�	ߊ���F"[����I�=�>N��ñn8�������4��ś����l�4�S��7n�� �����ݯ]�,;���>�7}�W������z7hO�����Fu�r_������'7���y�����,��.q�Ď2
����v��Lo�@CnO������*}	dD��l�X�[�,VOH����)g֖�?�jVQ�uR�mȖ� �*se�\b.�[E��	�8zM"�P���%��L��2�T	m�S�eb:})���q�Z����/ZӚ���9��
tpn���Q��6*��ɎL�3f��
���hE�24�LNH�Q�$ @>=�f��U�K��g6�}ie���+�FxA�uz�K/騡�k#ٚ҅M's��0�ё&iOM��I�������\�M>}�۶�9������l�;�jQڴނ��̊�>� 췌�`f��3���)�V�p��� +AY�O��W^��2�jDD�p(U�0Sm�I�x���s���T��0���06��?rJe_�C�'��c��	��6m�5<���PY<%�\Nt	,�i�*��قRθ���aa��#����8ňS�r����~���Z����<�n��\Z��}�Bu���(���a���E�D,���������H��o�>* ]Bf ��柎x�v�3f�7��WJ7B�:�	�\�I�kVG��|j#33j���\-�ڧY����S�\�{���'m���"��i�#��KK�Ӑt}�7��}t�D6꒥�ޟ�˔���Y��G�b��h���=�qq�J����I��/AҨ�����:�	����b%��|ı�%H)�އ��~�tn��.3�N��J��K�%v�H��%<~I��b<�m�9��R�QY�L�n���s�^M���w�&��D�iQ����$+�����wK��=D��y�Z^s�K�tU���@��Ļ��D�Rq����-6���4��A�3V�*��9"����K��Xl�W+4P��m�Y��aT��E��C��}��$�f��S���&B����)�D����X�C�Ҙ.�\Q�̸�ϥ�? 6�����Fʘk�ZtOu��Xy�Ɉߎ�ڠb�w��l�G�Q%.�eF޺%df���q͒��5��Z SB<M˷!^���:���ԥ����Hm�71[�_�)J�A��Nb�.�TV���-�؝����Y#U�C�\D��L�V��kG3�AG�B�dż�f9�O:u���cQ��'l�Cܨ7]I��V��y�F2���Qv�D��}E]���e�l�DK����W�w����(Hv�4WyɆFq�~�]$��F�\� �*��k���d��ޣw-��?�c�V�
yBĀ���S�h+<���R��md���Y�犽(GvO5NVg���Q�����Zf�0���&�o�F`H���AQm�_E��#r�J$A�r��褩♄Ӹ��đד���X�F�9���U���,�����ۓoY���p��A+�Nr��Ǒ���JM%��:�2��2�&�;�/g�j�߈͌��+H�0���_���+2W��k0��5du�Y]���t��u�f[4~�9�i.����3��,�2;�8���V�P�-��*�5��ޣ-��Kv��X
w��H'h�$�[NQJ��7����J��v�f�ӊ�U�~�
�3�j���?La��i	�:�v;&����S7�@8��U��g��&�g\HC�O��,��C�ΙH��DӜ�I�]<��}b��=�L�2д�����#�Mx	��ʔ���@�� ��Q0i��o�_]��2@+���W����wh����V��b�.�*p#F�T�
1�V��v���6lgn��"���S��ҹ�^����2��H����Q�Qa%KF��-ky�ݷ���T�GPB�>��Ζ�In=x�H�S��2f��MR���W���]��.y��� �wTvM�#��j2=͛2R�-�!$
��Qp�"��8l�B�܆��3ׇ�D#��K������gg>Y��C˛C^LɎ���/���俞���W�p̋qQ��m��b���u���AyW��y�ޒ(��W�1'd���7�zu:���#����vO�=\��,�i��M���=�@ѐ�K�Z!�w�[�_��}��VGЗr��U�!U�\̍��	��f }q��B�rUF)-.MAǲ�� �}(Ű�ed��2(�Ǘ��	��t���%SQ��}�drw��x�'�W���5#�&����*��ч��9�2ښ�����d��G7m6�9�0�=�^ V���c$�J�A�8�e�2H�g���%�s�5V_�w��!��)�C�Axլ�2���b�6�:�6N� %�߲Mbu��O��7��������U����crWk��R<M�����ٌmyl���kЇ.*¯��hߩ:�����PdւD^^t��}\����/��\��s����LLz�c:�p_��[�*������n9l��V��0����Xj,�n�*��%�kd�5	Cm&�si-��}��CV�*͚���/,�+y��pQ�wq��GY<ԏ~Ӭ^�o/:�po��t �"6��r�p^�-�^���ԇ)� c�i�T�����Qb2� ��[!v8���(�����R����&F ��s�m^I��R�~����`BF�{،zU����h�r�|KU�k÷�)���m���A,��ڥ�J^)J����Ӡqo��&�h$��ːt%*sw%����1'P�5�E��K��[�@ү�ۿ���e�e܆r�KJ�� >"��I�\M�P�E�E�K�VC7�,���K���
�n�?��� vI$�B��q���k9����z��K2/")q��#� � ��XȆ�Wۺ��i=ɉV�X[h�&�Q'�T��ԋ�V�!�ǅ(�GNl-��`���W�ʿ-�.Џ�kl�I/,r�A�@��(�G�g���8Ǽ񔸓�[�ù�'=�Z"��a2j�Qj)��=�TJ��N��Ʊ$6{@��f�;��Φ�!7V>� X(=~2��͉�s�7�!�����k����G�<*�����Q���FK�변���"���t�'T�L�S[[�v�kTB;R�T`1��o�:ܚ[�[�ۼd�g���!�$�(����6� �>4s���MaӶś��^s��QϾ=�u�% x�8u�#k�CN�΍Lx��?UD�)��,�e;��	�!�B�
�CC�~s]��f�>.�R�|ĥ����K�ye�m�8 �ߪ�I�m%����@�(�I���JX��.�.P��&a,�*#�i(�����������3h�e�ybzeFǉϻƢ��0R�1�䚣 � �˜��P��=CEQ?R(;\�өxx��C(��-�O�IM��d�瑡��D �R��pH�NλzeW���ú�Ae�m��,;oS��/} ��('����8�����\�\G�ަ#�,�'p��J��	�C�C��]8�4Ϫidn1Bgh�x�����%�.5��Q�,�\��vԵ>�r�^�`兇���;|�5�*hٙ���	�vM~~�B�"Yp�2���o`lإ��@t��T�_�ӛ#�n�R�
�	cڃ�TgG���[1�J3�y �y�����l���WѨ�`l�j���II!$�[�䔶(*9w��;�����֠�:��i���ί_�F`9�9��2Q�/�</gɼm��}2�G�a�J��oZ�Ø�j�Joq��v�wP����9�,���G/�]ݑP�\x����D��� i�eE�K=�l���4W�XŒ~[P4��s}�>�*\)��D�.�_�t�s!���O�W����1]'xٕpP¶���FE�.��)��� ��G����]�c\�3A9�*%J����8o����xKV���ɮy�����Ux%��w��b��U]�a����
�t�K��ޒ$0!�(����w�Ϡ�y3JG�ѿ��$��$�7V\�Q��_�
��\�H �A�>;���L��	Q�֤d�sm\�2�FVa�Pý�[-�n���eX�3�eX�ɤ���Hx��N%�d�|Ӗ����oPDx�
HrY��k
i��&���}�����7[�{\����n������(��A����+�`�D����k��˱�+�߶��d���D ͷ�MH�ۇA��`��F�^	aP��~I�1�
��)+��8<�V@�5�~�K�H�J�`�5�7��N�܊�b�=� �rC�-�(��B`a9ӦL�٬�t�1�5y
A2WW��n�~�v�ȬdZDm�z�u
�����n]a5�c�϶���)�/�\��g��N���z;��k��gD~��$���{����T_j�������V��%᲋N~q����(b�l��J=x�kq�Lc��/D����绠�(T�� -�%
�CA�Z�W�8�BF(���w����mxuMN�}���٥>b�����&�d3^@���V~��YR�w�J��`�2�z{��:�uϹ�*49]����\>+` ��r�T�h�:x����T� &zz�✗�d�a	�ʑ�����jY������tÊ?�c������� �+��+t2*[#_�;%LƊX�f.͊t���Nw5������&E�70Di��@�iTq�����e=In�G6�`�r2�#n��f�
7E�ғ�=������5���ׯ�0�����^�����M{��g[ŉ�=�F
ݼ�"V���:��j�
��Z�!�&$�3��ߋ�u���Y��\'�,T{̞*��b����f�|)������� ��K�~`��~#Q�F}��7�x˗��e���KH�<ІM�^�\��6����I2�L3��C�b�h?\� ����=s���i�0�!��E����-n�?Ō�6��f�S�Y�PM��,����Gj]�幍@ �ad'�@����:|)�`WG:rv	S�f�&�t��VQ
��YV����|*M����ნyv.Oi����>Y/��gS�J�}>�LH��@$��|!�)|�1�x��Q��Fb߷�*�m���VvƟ�Ǜ�oꚎ�שHH��Ϲ~\S轱�J��͔���^ v�F��:��Wl���t\5�E��<֜�h��MJa��.v$` ��9 ��	�WB�b�+�X|&�{�F�`����4��	�z��s����d;�+�xk���F���!���{�k8�[ɑ�:���%o�Z#���Y��m -���L��X%	T{iɞ_$x��ѫ��4S����÷� g'%�l<
�1C9Z`�c�����k��q�$W����@s����v�][��d����S���05��������1����p�l����/�M3�N3�����߄���Zc"�a��!�BR�0{��J�"w�O&l��⹥�3�.��hJ�-�4f)�⧍9ޟc$Œ���ҙ=[���0�&�Gj$�r #X����B^��ҘjT��J_i���_�c[�7�X��'�9I^U��1�w�Ԓ��z=-�z�3'�y�w����R;�֪�����%�F/�V��O�?�|�6yV]��V(v`���{��b1d��H��0̂C\q �T��]�	�j7E���PǏ0�Rp4��������sdz;��Z��N�;�I��J�D�	cJ�L#sYz*�@��ǓI���ɜ�_��;1ƧYd�*��jC��e�]�/�FQ���K�b?�f��4�K'�iDi e�T��hG!�[��‽�?��3:+{��>{U,{^��mq�v�KGr���eVL{�������#0�  O'̉�Cz�,e��B��8�@=]��?��o�� :�����Q� <cˑ��	7XE�!�Y�~d��),��ه� ��������Y�Vo.a4f��=��#��C��GV��I�
k�YR&�V> L>��4W��`�`
��68��%�xJ�58�wk���z�G]���a��J-���앍�w<0 l����@�ό�f$����'�� O�G)�*�k� f�KZ@o��6���Dc��.�1",�ZK򂋫\�[M�!p�4��%`���N��q�$���ǝ� ��<%�pvO�̐å����g I7��C�gL���Q�r�T�����AX`s���-"�t��_uT퀏V��3��	�\�O�`t�U�q�|C�H��[�-�s����N�"�0��� Nn�X�t��*��]��G��6�Y�<�%<���O�Z��r+��� ��#��@�5B�XC:�p���q�oY*M3-v��b#*��b[lXz�Ip���P\�e�2b����CUފ�]��v�Xy��JH@I�˥t�[��p��ŶKP�9��2��6i$t��W�Kj�Vu��b2�l��5�Le���Y�r|kP*՞���E!׊ �d�����W�dn��������a��UJ��S�\NƸ��G��=^W�Hw��}$�VJ C����/ۂ��xa��1�{����mȗg�K�V�'�=�O<����ZrW-���1�m��zos�f���3��f���t3��������-+9t��+�i
�c츳'CSo�:1�{�,�1a	�>��[�0��=�IE�>�yo�p�^��!}a�ߛ!̯9��P��~?��YZ��QEAl�+�s���^�=�w8\ɫ+����F����<�����8��D$LB����E�	��\���n�Y��/B�R'��:8h�l�<�6X�S$ d
?z6���8���hr��1�@�?NÔR�M�T�����|�����|S�Q�k�A7��52�ƺ����M}F��Tb�ʚ���l�;-e�e���WF�Y5�3u��y|<\w��q�A'�����Lc��jF5o��ka�;�V4AT���)]�$��<�*��g"ჽ�vW�8Y3���	|?��������>��^Ɨ���4����l�v��jB�(�Yzf�n��0މY�X����аH$u�<V_̓�@\�x8E
C����`�nN��M�������7E��߫	�F��RZ�ڠ�� ��hi�����o�'�ݳ^v���+a�C��U�R�L����3�O��m矺�(�f.��3�!��z��U:6Xw��`�ϘC�����՟r�
�a����G�P%��j��"H���VΉ�O�_�k}���ϓ��GD�V϶�4���Gr1�	}�]ʬ?y r��Y�]�贤J��E�^��T�������ū
��-�a����H��p��g3�N?���ĤJ��/�m�!$ 1��[�l�ȿ���y�����L��� ��<��.�W�B�Z���6/������y�4�jb*�ꏞ+`��&�3zFA��C��~\׶�0a�����ZhĴ��0�v�l�M�D�爖�o�t<5�ܝʂϗ�,z���ލ�G��$D~����I�d[�6�j"����* :H��Y�
U5k�h΀^��&����Y�F��[-��°v�MJ�=41��K^y�dj��:gm	�sH˓�L����F�vv=�����gp  �Tcj�k�o���}n�Ā��ǅ���&�|bz��Ӟ|�������,�Tӎf�A{Й8�*j���M���.�E����X�.��i�i�we���~S��`QB�K(�^\ad��ΓN.�,�9���Y����l%`�-%8��˒�`�cQ���XT]�\����)�0zhi����쓔����M�<�k/iuw��v+�jٕ�An�#�\�D�!Ma�#���v� V<�hw{'��b���m� ~\B��&1�A���韻O�����)e��l�al��v�%;����N����,	���,��I&n�?����J��wC���B}f<�ԅNԈ����ƞ�1���;�{%���[Y���uTt����9���P�����E�{ۅ/(�0�V�d��#��[~{IL=J2b�B�pm�t�������rwcsl��T�(Xm�L�3\�ČFZl�ӏ��N�p�;9���C�y.B9�mRp�����*8�<Z�ѱy/pǪ�P�6�Ba)����Da�s�V��k��`�y����M�b�轿��")�f�t��~,p���'�M�3M�P�6,4�=�󱅍�m�F֎�qq�!��Z��(��f�e��̺��/�NF�CQ�f��b��|ǟc�1�������j��l����?u�e,=��`�Sߏ7\/6��B��`F:1
i����71���Ъ�N�@�)`��H
V�,M�E�'�ޝgz4*�_��ߜ��������V�^9�3��H�
����F�W��g㔰�.��}?���vz�lȔ��A$����܅8�h��I�y��~F)����8{�;��=�c[��i��T�*8�L\�h�w�|����e��w3#�͓�7�G���~��!�PI��T��b���V:]�/���HU`+��\"��@��ZK�F_c�M�q	j��ǲ�����	H�*�^h�n��U�K�s��So�Y!���V��8��x��M�2� 0��bP�4�y�[k���pq��b��̳��$"�@9CT+c�Q��q�i�+�7����"D�ޫ�_��,�X6��XG�� ��㠷;r�%����A{	����-��,���i�\��(4`�������E�a˳��"���7/���X�v���n��-�c��!�3�v���hW�ӡ3L"p���83�57g�(o�ڕ��J��R���B��͟ χO�%�_����@|��T^������*�!ɥ͟c�3R�~@^XMRM�Y�x�zL��>��O�6vs�R���-,\@�'\3@��$Ձ�Q�ݬ���������ı��g��/��H?=[4�k����]�;^���g���5��&S̩h����]j�;�J2���N;��w��ս�m�]�Z۽Ln�`r�{twz��v�h*��@�G!A�݆� q $GrC� f�VOƂ�Ʋ�)u�)M΁����F���`�2���揬�xv��.����� �w.H8e|x�C6�x���:G��3�.� ����%������ !��n�r��j���Z�����4	ga�ؐ�!���7��Nq��Xyn�Ö�@��	��ب����� ���s���JkZ{'��)T��*��#��z�O6�j~�\�-�u���1l���2�_b_ȝ|��o)��ܧb]H���U�6J��Q^���L�E1:�k��!����"Vt`BU�Pŗ�J��}(�r=v[*��]��
Dˈj��i����N�qP�lMy�W}L-��P�BN@�q��S�,[*��1�u�ӏ'�C�������>惣~�,8+�oi��;���8�#�? �<|�xך�+?��VAu}.��-��w�z��l�8V��^��,_�9EӋ��x#:Nĵ�Z��x�8��ue��W%:�kB�F�Tu��U1��u�Y�4�����u!�4�s�G8gê�:˞>���\r뫖�@����Ju�X��C±=6��У%�l��D ~-��F+�K��6=ZR����4-O�,�7�ֆ֣z���B'Z�ђzρ�4����r�y8sg.����,T�h)��V(ں�f����ߊ`}�J���vћ��y^��S����� ������{�*e9��F�D���`/y+���vO, n���g��E ����!\�̳�|���6��lr �ө*jVz��6ض��}Jt�w�s�G��I� ���64y���``��z֩K*k7F��������b`/)�^�2�^{� ���|��V�Ѧ*4��B����ȱj�+n��̺�������38ۜ� �.��2L�9����L�07{K�}���>�6N�$�/�!�[~�F��_XhK ���Mi-�ጾ����6�3kN��Um��\�E8 J�'_���O9��w���i��F
w�6�!X7��+S�h$�;ü��'t�|w`^�B&LD0\�$�n��$�@^%����̰t�Ƕ��1���h>>�&���n��Ȥ��O�BU'+]���G�k��K�xZ�Ĳ����`v42����in�̙A;�F���tj�`s��i��K� ���B4.����j�^_o�C2~6�����,���	��ٹ�L{�4�ľ[������n�^kO{{�،�'dq�m�7�⨿�.0�B|�a�"o�տ̣=x5�+��:�Dt��
���*���|`��Z�|췚_�56�� O	B,�P�aߕD�B���@Q\���n4aJ���|e<��^"����̲x,�������������{D��Z�g�y�io��P �6�"��y�*"��m�"E�x��:�!=�V`�s��oʃq��81�>�q~;苞��ϻ��0H!Y`VD��~XF��=�{`�Ɏ$`�X��<��P&��
��r�y[�gx��,=�����N�9��Ep������_^B�f�%�4,W�&��{�b�˿Vق����?ϑ�;�����,�Q�)hb�=䍛m5
�>/�{U~�RQ�5���s�e�*������,4��f�Cݐѿ�I��p�{��B�ܔ[��:�	�(fm	{�������>	ˌ;u�^������w����p�$j#:�g�l8=^
�^���ȉ~��+��#1���ꦉq�&�6&����-jf���ث.�l�}�
l~��`���;�z^��yY�����\�7	����Xb��`�>�����z���]C��FPc3��o���~β����ca���3uM-H�U�e�uy�?$\Ǐ����K�� ��چ�a�>~���j��'6pieaQIL�w��*� fcB�I����1h��I<R�Xu����g�*P�$���ۯ�;݊����I�F�W�M�r&�ș��>/{"�#uJZ�vB���;��wG�c���q���Rw�VAB\�U�x�=��5�y՛Q�m��,��.���΃���i|Sr�=v�}��w �<(N-���1��!�UN:���Xd�{o���;n|�I��Vk!<�<�1+{:������k�?���|X;c#��ޛ&m�ښ��JT'���_�m��8��Oc����%��Jy�<jT+�ՠM��4�C�}�I�s�䐧���ˢ�X��J	2k�W��*��z?�s�~@5���;�)��gj�?����oX�wǣ>ʰF���+ͶLU,ڎ3b�(HϤ��������������uw��?ZC����1[�
�
��[�Ήx-��7Hpq�ߔ/Mqjcȷ�G��iM�uo�~}B\ `3�?���h�HD��kI�_�c��"�ܣ��R4]/3H��Z'+�|��}E������a�?٤.��
J�N�rq�"�S�]-}DU�Լ�z�%���'z�[�Ҟ�Gl�qA큨5���|�\F#����j��6Њf.�>�!T����B�\�?_۫�U�L��K�[sev�� 3�Nwo8>�x��j
���E���/Ef�(�� 
lC�ơ8/�;��-��S�O���K^��B�b�v���b���A��� E���w#��9}�C�}��|$�m�� :�Ճ4'�>�ĸ���j��uc������T��T��s4aj��&v7�G6��:ϒΙ�k�*�k��R
��ș�;I�����{5�9)ŗ�;����{J�W(1[@���Q��1��(��)���9���&x�r0�o(���{�=z������&�^!S�8�a���A>�]ے��4D�'}x}i��&���8̀c�@�l_��/��GL����V�[]����H��>r��1	"@�5��@$U@r���0k����RZ��o�#����+�a�"@���R��}!# � nP�d�؝E0ҷ.��G��1����\˒V^�BS�͘��%�_j�ɼV!��>2��:0з��g��H���^V�{Wr�@Ů���A~���;R{����D�r�8tY�~��N|�F���G�� ��|��1]xU?�iF�����`��b�m�ENh��J�����}O5Q��CŤ06��$i��J�`Ǖq��[��4pv���ɬ�� �����ׂ�����鈯,e���R؜>����ֱɭ���a�2,R�t��8z���럟���l���� �4#esA��P��}��O��4|���](�^��Յ�?p��L�� d�kl���_Q	KA坐�Y|���C�/D�"t��B�[k���8h��&���f�F�d�Yxk%P���Y�oUB�����ˤd�����������ѷ�*�F��L�>�R�|����M}��Lz���{� ��:Q�0^�S��5tGk	a�a�mNCL�p�L"vˠO}w=8��m�t_+j�㯒O[�YlZ�7�%3�PN���V�T�T���ն^.!d��#�|G�,�}��R/��i�QI�\?��Iv�.P
3�Q��6+`<P�#�qk
ӯD����L�Ȭ���-����8S�OH��6
�pN��TvJ4���;��;9:�s'�49?����+xՍ���{��we������B%�]I��id4Y[�h�u��������W�|��O��ir$��K+�z[��#7Z*���{e\lM׎�D��fPH1���d�iR�w��*~h|-����i�<�|��+��=��>�(���o�#����邑s
�h]��NO��1��+s�9¤�b&��j(w(}��t��e��koY;1��1m���G��/m�q� �xf�_�D��ZS�� XW$w�<6Ui��e�<���`Y�ݙ�P*�+p��,��̚9�6��_��%tM��ی�G�Vj����� 3
;�ܿx���}�4�@�^�0��_>��o���i������FS/��GޗD^��=1T�
������[��o���q2}�%�w��b���Ƃ�9�ڜ�|wwMH��c;s,Ć]5:�er;y1ɗ
�%�^�\᣼<Ny�s�m��L�nT.waMѩ�z��j,H�M�tZ(0�c���Q���>�uݖ�S)t�b�/PY�1���n簶P���L���b�����˩ͽ5��\T���~uP�6�	Z��0�f}>Ls�c�2v-˾��ఒ�%7�@m'���	��SW�.G�x�o	����1S%�,�h�e�~�8�}cK��&���@v�m��*`b�M�k�6�.���?֎��aF�Q3I[Ҽ������/�Snd�+S6�����9LLD������=Я����֌���e�W~ߒ�Sk�X�Z�=�w������;��d���K�h���G�|沏���_1g�R:�ga�p?��Η0Tqu0(8[@^&��>��2�i����.Lx�H����(,�W7�i��7�|�(����%����!���RЂ��7��^8l�����dŏ�D�=��K��:�V��J])tI<���m��PS���s�����S�E�1�Ն��Lbf�>�ѭZB�^<ڙ�X����"m69�u2�G��gc�4�X`����q���c�:Rk�z���/v�
��v��X����w��]T{j*�O�=�ZGEk������g=�x̍թ�3������q��.�6��(�ge�K��L������P�W��<����F40�`�s:Mx�p";A��4����ա9��Z2>G+X�|��1uݥg�U�\�^���}g�"Û��9PHo�<�Pn����M����6���&�<~�˴�aw��?1��$�'�j#�f��+�	a)�؊<�ޓod�0>��p�Lh���K�w�J�"�.�	��Y1,���/ot��i�����kl��MZ(��p�i$@G�p2�����]��I�{(-/
���U%\s��xbx�Wn�$z\��y�E)��
�QYk��X��1��� q$oy��-rk'�����x��3�S
r��b�|�!�r7nC���&J9y�I�)eޞ�֝yg�����(�GwOՕ]�8E�COu����)�JZ�,X���V��S�U
�������\϶��2�5�Ep�mK�ӗ$O-6��|���r�/���W��i���I����˨4����*sI��������
�h��/��֎u��հ|�b��}s?iEJ�����Ġ�.���4g�ҏ~D��y���[X8�O�A޸�Ϗy�:w��}}����L���|ya�Q�&��h�e����񏭏�Ĭx(P�};=7-��L�C��0��Tk��DL�!�=�E���7�G�MPX9K����'�b�O��.���g�4*�8�	�Ez)���R����Rε���ՒI����
��"c��B�q�"
��g�捈:}�HNT��>��A��#�#8ɏ��d'�Z�hN��m���XUF�ɉ~��n���S�f��j- !�@Q���@T�dA ɭ7��	;�-խ<�l��Z�{_ ���Y��Gb'�jP��Go6V��Ҽ�UY�jJO��4�����F��2��Y7��*E��q=�a);��]�]�3�*ɦ`EXb�8�q���M�FRX�?�Ɠ ڋ�P�=��M�%uu�M���\)��|�:LuD�h��7����c;[n|�����sYS'�Ν���b�D���i���[*��`\�Z*�z����<��9}f���(tΐ|F�C$ ���R��qA�:X=#�I>h�����!-f�æ�*��c�-S9'm��6��b��D?���!y�$�Q3 ���pJg���x��M�C'���]��A{� *��{�8��(�Yd�'!��$C�&��0���$I-(���[�ѧ6� �%�/^��$c��� ��@�)��0P ��(:)^|C��d,�M�ik�7��y�\˻ ��'��R-�YLcP4��oc��t��C�iɴl�k��C��2�u�����a(��)�fL-�]���}�����if4��)�@���[	{�p�������x���� ������קʾQ5`i��X�(ߤ�&�T�©�O:�f�p�)9��@Jc�W�՞c��R�~z�!��M�5��e����Lg�QJ�����L����3[�G�/?(	�޽�d���eR����<?���5��:䄨w��@�.Ե[j3��z$�l}lǮ8��j"��!}S�T��	����FSP�c��GH�qc�i����1T\m2K�T\�WER��[Hb{�����;@/n�|��b01��X#G��cJ��d���ciUDn ��7cI �G齒�*�Fè�Β���NrF��@���]�P���ԑTu1_I��g��H�Ҫ���W˱@��Z@��j���䈐��M�H$�0X߁�?>Ey�ʡ��}�5��'�j��TY�h�CJ���[��%�z��/n��ZA��I�u��ej	$�+�)4�!��ك�o�hpKf���ԒݛrI�~B������F̹dth��e��qi?	�h�j_,y�Ae0L�7c���f9����X!�����!`�@����K�>�r���]+ѹ���s�Vv���W�}:R�> �?��@gջN�o0�%�*����5��{V�r�~.>��smR���.�P�
L��{�b���ț�%j����C�Qj�C�@�v�~�X���9�:)��Fk�{v��'0�)���1��I�Z�q�L����Dv���r68:���K)�6�9��1���t.Qj��H�����=6ne/���H�6��n#>�-�Z�V������w|�!�שϝ�>U*��W./�����C�#7g:�l݅��>g�<�f��9U	�$U�%ޱ��~f|D���Zw�wY7ʜ~��۰��%q����2"��,x������9��V;�FǼ�h(Ĺ(;kӝ�@�߇J�:p�J槴[q*kPr� n���;@ԂS��3I���>4�n���W,����h�ƤKqV�g����,� 5�!��j���A1�Q��}o�:�,��v�d�vs�(�Pia<UF�^� l�U��)	ٝ�Ql�� ���v�j�\�o?��p����@q'���
�F��r��Qq���E`�lG�&V�2N�I>�o ���\C��؜TB�zj�Q��"����0�U��ؑ	� sM��V"M�:C�Q����j*�f�c$��
>��B�n�����tL�@U�)b��|?O�xяy]x���e[5�u¾�]����P�U���t~ia���!� {7:��N8xVS��:�ם��YLZ[nĕ��NF@�`3�Ff��V����t� ��D�)�f��7���[����AES���+ڦ:lW���CN���]/�9/��q �*(?j�Lc*Wϫ��)c���Ѻ��y5��?=V?���<�k�M��A5d��A���y T�BD�� Z�~��/��4[7���^�>��>�݄?ӵ{��0��o5��vU��bFڔ;@�=�S(�n&���*Q5��MrBb�V�Q̶�N���рITvZ+�y�X�f�I �a+=f����,T�)<��e�ؽ���f�c3 c8/[�T�������Λ�E��@Y�����p��� Q�,p�&��sl�\��L����uW��s�'�B��jSq0USI�19��靯��5-/�M43Ʌ$�X��&�U�J???�֓�kE$��}�5���Q��#���@<�z��<����[O*~|��r	�f��1<� F���]��;���$�c{���sH�˲�v�	U��*�E~�WԱ����#iS.Xݡm�5�7�S�l��Z�:@a#ܮ��@	l���&�o���c���i����,�we�S�8���ډ����tT���j�Ȕ�UKq�O��O���8��#��������x���"�6���lK��&�G1����6R�@}��,A��/]�0j��U���=�O˩�GӇ�/�1��t9%`�siw����q�ݲ-��A�5J� ��c���D��|!�Ľ?oα1*$�s{�:�*b��V�JV	��Q�u5��`^�`�{��ܧ ��V�m9����`g���JE�����n���<^�P�
�
��F�:��.�������p�� �u��M\�T���٨L����L�P�u��8�iiEK���ʑ-�Ml|Zպ�r\��֙���^%qC>w�0w�q������
=���N�[��l������tsI(3��aJD�N�����ci`��/v�Rh(c�J)EN�[i�/�[f'pD��,?�"�
k��0>	ʄ�Z0]���o���_��������BU�2�d+���Z��;�2W>� �'*�TY?���h>�'�?t��� w1�!�_�ha1�(���[�+��xF��ޱHx��a�TnRC�İ(7t�Ȼ�����q���;3(�5>V��>Jˤp�t\�֝�|{۲R����#��t�S
�����wz^�wj���&@G�KQ��z���"�0j��<��+��d�I�.ѩ�C������-K�DX��I�`�V�F|����*_{�G/Xݤ4������������ i~�Fb���SQ�-�~��h�Ek�����.�����n����#xH�Ae�f�O�EAy�d7*((#�VD�n��N�J��/�������L����[tfi�a�ORN�`cZL�=[�#� ��8n\˳��ca)��y���0:�[Q�wu��v�O2z;�d��c[��W��rF��p�.F�A�cֆ>�~)��~���ƈ����<̐N�MM�A:���٣�
���j2���w�\�|��c7�H ��C3�ClB^�چ;�IQH�X� yT�b�Q�`z'�@��lU���ox�qfꝠ�0(l�/�-~}��-�f����e��dP�g�?	�VHSXjh.ΘZ{L�
l:�맧.��,F�v�w�`C~�H$�Bp���.0��xdi@8*G�R�G5�E�^����� �� v=)]�p}c��b��JL�=���'�[�3��R2$ZT�9�\����(}o�]����X)l����Ϙ�j�&���ܡTs��.�ʸ�Rʦ��z{I��~nIB2�4ߔ�e���Q��R�/�e� �IBZ���=��	����b�[:�)$^ �Q���~�1%��o�5n�[3��D���`䝏�f�%�2�7�fp�9��bP����r�*"�~��l�!���-�Q$�O��+�S�(z��������Cə�  �o~�G�@���s�"�m���S���,�>7��(hǘ�'�B����@�ʊ^�F��ZJ�u��{=ɪ���6-#���8�:���<|t�����d�s�F����	���W���9(v"���H.�Gz��`|$�( !����eDy�:��� zɞ�IӺ�+���-[i�Y���Tb#P�e �,��n�Q��������<[��lg;��~]�W�0��0�&�'4^s�H���A�}v��&ݒ]o��]Nˣa�e�~3v@�P=�J~�x{�Bcْ�҇2427'&������f�R��ک�R!��͉8�=��$��M��߯\,F���x9�2�kl�������kC�
&�v�=Q��KA����dP����2��`��a݆~�k|��)�H�������ӡP⨞���Yg7��jƚ���t{gM��e����ф�5K���)%RC����*=g�I&���	�g�rک�� <}��Ea+�*��#���`�?��،[��z\��䑿:�'�V,�.azqބ���h������xJ� ܶ)I--�O��vBG#�y���z4��#_J�൚�<�ᐠ�&��0�$f�D�������i��ّ���8~v-�#[��������a��Z�y�)�a��7F߁Щlm���([�#U|��(wc����ŮF���5,�	_��9����E,�댍� qD��3g�	�E���phw��!X�ޕH�j�׫C����5_*���T�_�m���￣ �UJE��.�|�+0��[!+�w�+c��i�h���j�?����G�	Q��Ŭ^-MzKV��W|j;ڀ_�	E�$t�"a?;^�w��:pנ��l���.�� I[�#ujVX�9.Mqu5d�Vy �����^aҺ!��F�|��.�BhA�6F*QؤH䏦Ĭ��4�U��I%t�Hu�����ҤXe���Z��.x�yd�P\+�:iO1��#UH�Sj��ӲQ�x7����:v�k�D�����Z�C���+tǚ���e(�
��N��6��3��YC���
�tK@�˹��"��<l���S���%���~��
�^(ϖQ^OT�˛pP�(��MMu�7����3�B�\��m*�����,�
�6f{O����:꥟S�%���2B�[���r�s/��hTG{�m�j����+Hx�@��m�/6�Qص�qL��R���a�_��%S�`p467&�SPL<Og��u��U(ٻ\Y���J6]�X_�	*O��_����,�����,~� >p�cE�����;y6͓[W�B0�~���bC&�ŕG;��$:�@�':�������D����
v:��p��Q�K$�������k�C�\�RE����y��OC��]͸Z�E����d)��E=��-J�w��S#��ə#�$����[�#�m��*��� �׸�jʍ�O7�%�G<�ߒ��'*�I�YuS�|�]f=��"o��P%Q�|� ���`����GRd� �h}g�����'ܧw���9tg	����O���:)�'��3r�ؗx��N���t�_��������Y��O���Z-�t;��� UhB�O?�S���VY��a:��p���	A��3����h3��s�D$ӧi��pR��1��#�H�d����B"�|[�Ô��w����V/F��zޢ|�T�8�X=��FϊI0~FA'gf����"��)G������C�v���H�d��2~��~�cڃo���i߾���=��x6``߿�[f�e��9�"�e`�"��ץbbK�`}�	�6����Y�:}\z�jF��)z�%v�e/�k��ù��5�afi��T�x`X�}p� nH��se�P�� g��MZk���`Xl# ����*��4z%F�W���M�N[+�4-Z�9\�����,p���=3��9�I1��6˶{��j%?�f�E��R�OƈC��z�[���{ğb�X���fXے�l+իfZ����sDo��uXv8qh}�����92k "�w���'`nM;�'�=S��R�i���Cw�2��F!�5d����.זu�o$-���m����&��,Bu���S47C�V�,�kӝ5	��j)<�6��|�:3�[��n��,�;\keV5_�.}�(.����I�gf������f]�R$Z���I�ۊˑC6ҷ���s�8�]����C�~Z0ҿ��=� �� b��=��9�&���> �Ub)�]B�{H�ct�&���'^Oc6[��7t��j���FX~/Dp`V�XƗ����v�l齢���Vv[hv@�+,v�\�<[�W��oG~�F�X��c�u��bKF���C��$��T�~~=��?����Ķ��n$����l"c��l�)�ĸ��������2��ǘx��y4�h뉈�!u�f?JR�'E�:���s�e�1�n��R>Fr�+C��X�4^�$n�)�T�����3�=�Co����@�V}IՉ{�� @1�'�o�d�EW��iI�Dp���S���)8UN�)���H��B��3Z�����s)?G�G���&?!�����CnN#�N�B�
Rќ����
�$\0��r!�)�t�A��+=�/p 9 �Y��Ӛ�V�d���M�]
�PL#�=nw�@&�֍���=]7�3n��~&�����q�����sE|*����q�G��)�w��R$��EQ�u�P�/��U�hSj��21z�sl����y+�.����9��CO����=F�6��k��;���a������C��xeZS *'�qV܍���cm-8�<�����4�"*�z[�ǁ��;���a��+ɳ����y�ąO{��[� 1�\/�V��ܮx���7�L�OH�͑Wx���P���4:���.���cU�]���7f��o��ӯO/W�|����Gqj�q���e�Q����e.������^���R"4c����>��_O;2��%^�Tc� e�_i`�H����/��c����������Rı?�m�X��m+�S�0�X���ꁆ|e�h���-��jެ@"`��WK%
=Sb,Uj�~�%	=7z�����/^�d�@V�a��0{~⟘�"��i�In��\"؞�-a�YnA9��ά�pHDٖo΃��g�=�{yn��T��������W�$������م�����F<����:�F�z��O]�v�
2�D$�b�R��f�N �џ�4�P�<q||6�!5��h�))%�6��Os���� ���j���;efZM1@�L{S%�^��� ���Q���CP��tf�\cWsuq���Zt�N���:A�C���8��繅%jg��j��4���"FK�d�fb=���D���$hd�����_E�Yb���EK��@�{�����&�T=�������9��)p��j�����3%���j��(�U�ˀ|F�ւ�4O7�\�S�\�h$5у�?P>u���c�&��-k�����X&L,?d�lG[�F=�i��,>�?t�ۛa��a/\i�9ᆷ=��̟�Sf'w�9:7M8铁&�vJ#ƴ��rʎ�7!����Y�bGu�������%[�r�V��Sv̄kؖҨA.F����SqH�ɴ6B�K�q5Y�II	��$뇘���������S2�j��R,��D�����E�����_�д�V1��V����aOC�׆b�g�+)޹��4�>Pe�{~%�DH���Җ��בmi%��(�6�\��$2���w�|��/����F��B�M�;�dKZ_�д��ez���C����wN�Q�І2���
��)���y6�O��v�s�n^��o��6�/�_ͮ��s�����p.�U{Ć3G��
�p�]�jk���Y'�|=߽'Ε�{�-~��D�:KjӜ��L+~���#rf�Ҟ�z��q�{Q�H���f�zpWY�i��l$g��3~` +��o���b�LaQ�q�1Q-���4�]�(�+ȃ�у\�O���D-�I�**���r��;s~��@hx˞���6��실U*^���^E�xD������	�d.[�=f.7����OR�*��j��_w-�W������8�P7���7�U>f����x-:�-\��~��"�·@�|�h�S��]�-9�0�qZ:�y���d!�~��T��d�0�'�i�۲�Z��6�\?8\�KF�5�8��$`Y��2#���-kq����
5*Y���)��Se�-�mq���|�J��y{d���ue|��ڹ���߼>>�<ދ+S,��Z�\%l~Y�_#~�=�1q!���92D��U+
�ť��c=���ޒ��#6s��ST���5�\�.�ĩ�F�/��Ao�
̬e��gFy�}ڨ��zO@�P�H��-G�3FeN�S�Yi���{��R� �����Z��Ϳ���6"_�R��_n�3S~��xR�1��r�C�GaЈ4��
X�CB� �񪗈��=���8�'Jt�c����B�j/�J_x���mPoD��h�`�T��3�æ����F����+���(h2:QU6����6��#kQ���!�m��BP�L4���(�\��]�� [���҆n	J^�	��Q�������l�JR����ij��[�]�i䉸\Q�4�%�x�dӎ닰;�&vX,��m���Iﺛ�Z4�Ny�mq.���ﲤ��=�{o}T�m�iڹA����{�%��Y�%�e�:ȓ��x	��Nb��2�vv�$���t�_���롞�ܯ�,��	G5J�В۳_�y�6�=�^�n�""�S��|&��B������5�3}� ��ʶ��?�Azw�V��� �H��{-3�ju�<$%�����˨a�%�lOx�(�褉�=���L,��� ɏ����.�\Hp`�,����y��Y����W��o:b��@��U܃��A"���q���4��]�]h*�M��ƶ>,�Z\_��C��ƥ���|�dus�n;Bs����]�2�%�jN�
�4�����2xA��OE�l�ϩ�5hx�e����^���f�S?�T^-S� �|��U�T��1��`ћlD�MQ	q^�f���=�p[�3%x�+�ZO�:=�&9<�6l������X�O�|а��[��2 ��fCS�n�lJy�O�BiI�z-���]�盆݉0H�v�;���r%�z���e�$��T���'j�I9�6�<&���D����إ��/���t�|T,iY�� �!�^�������H�DK�Usb}�T��5y����Gv܉�媓��W�A��j%��3�
L!�ReS(�����.
���"�΄�8��|1�ʭ������)�5cB�����-[����~Ԭ
���c���LB0FMM�m�Vmu��j���A^�f0���L��*�\F���N��a��F��p~l��j�3IT����^�?(�1�h� 
�i�A�Y�r�R��.�R�z�a�0%@����S	ǅѪi�(�In�t�v��;u6�yz�+����~�&�o+ٵ��n^����Ь]�:����_�fJb{�Xj8H���g��C�	1���"���ZF��?�a��t�j-_�u��Ax�ˑs��F��rM�����:�mW2���Զ��>�: r!!C���	��[�(���V�" �g.��D���d��fƩ*�<W�PYc n���0c�������k5�B�5EF�&�NU��CfW>Oc��<��P�<\�It~A��a�M_�J���@��A�T�U��!��?L^"��J�e���U�(��жr}6.�B�i�yi� �H9d�w����٣��dA��x8jDE�{9�O��ځ��t�K�P�a�1�B�	t@%4�%�ۅ�z��.�8Q\3T�v�x�>���ՕJ��'�)iI�K�)�
�vg?u&ggL�
6���IH��X�
e6ro��%�=^�� =��[
Z����C��r������s�~�|/�~������xڏ�,a�K^�1�Y�|�(��[ͭ,��N��l�����%��]��r6�2vD`IFb4������nO�Z�E�.�ӕW՝�¹N�� ��m�����G"�Eԯ�(ˇ%��}�K�DkQ������F��,+êXH@֖�����Y<��t�y=ՙ��u)�'B�
K�a���Z3�1���0�u�+�̺�{%�Z�`��j����^�!oZ(������y��F�|���UP�hq<��^*W��n߰l����K��'q����>�=v������� :%���{76�QA`(�X���Xi7ÿhb>��޾�Z�����U�غ�1~0B��x�Oi�y��y�4��U]�T��<;��2}hJ��\VN����D�p�g �O`q��������ʢ����U��i.��F�EK���4���RH<Z�)�In��
W�D�f���^�~�%ڶ����wk��T 6����G�w�^H�H�EǨA��H��|�� �K�Ez���$f�B��R��+��N�N��2�שqn����AF4m�^ i�ۓZ��c����x�I��.�%����i�fb�$B�Qcr�l�r��BZ�[��W��^d�<O`�	&�f3����[	�WD�ҙ���e��������MC2�*�$��/YO 	���g���� b��c��~���a��(����3�V�1��iD�;>߹���!�i>fj��g�� dCZii�e X��P
�s�Kx��U�⯓� _��d0�z:��<����D#]JP��u�C4�{�?7��׎�"��=uF��tbS3��)Ǳ��!�%)}y|w� �szݬ�N���0���o���Mƽ'��š����)�2�u�P���AH�_bY*��=A*PD1Rj�[���­�N�4#�ӭUPi�=:���Y�G�G@�p��d�ѐⲼ�8p��;е�D���Eba�8�F
;��X�/�[�l$�H�U��'�$�kJ��G��A��?b.�]�\���ސ ��z<�]���Ў����[G7�$�w̽��w�q�ɯ�\��l1X��n�"�4Ev}��Ov���{����ՙ<yO��C�E�c�N�K2nRnw0kfDg�ѳ1��)�����&��#�<su����)����Pg��9mO�<�ĥ$�r��A�sʂ;,�K�R�k #�"�e��j��lF��O��p'��h�*�hW�/�����}��@�L���q�/�T��� ���B���b�s�u����,"�tcm/��q\w4%y$�x�9g��+U'���aD�Ϯ�H����$f�L�1���<�<�R��hd{t<Ҁ�*���M���SH(Q/Sև�0�?�&�e����䐵粖��O�K*=a֎'߹D?�Ĭ���,�팾���!j�0o�P�e/~�O��5�Ɏ-��rg{�"�{&0c�z�ռs�RX��D���g�K�dL�"�J�yqu����sQ���q��h}���㓔u�Q����]U:���mqG_0Q���@��;�D����{�-̀���\h�o�u��Ұ,G86c�b�X�+�rK�b~s�'��')��M]�Yڼ �����^��9S0q�Z���R�VTV���=��R`�2I�g>̃@j��ׄ���_��d�9)���wQ�h���#e���*g���x�nz�����+$7?���|C�cLi��n��"��k:��J���b��Y�I�]k?Lba[dD~K�1��Py��"p�$%��fj�A����7~����cTx��p�㴼�m������詧96������y��体9S��L6sk$���צI�xA0�cςC
-�[%svx��~�G���#k�|O>T1Hя�fR�D�TV0"X(�R��Y�<@��F���u�K��O�~,/���$I�Ⱦ���&�Y�l�Yͼ�|Ω���]�f��y��:�<B��̰�b�	�k�0�T�!� ���4���l�I�ƞ�N9�7�b&�>&}����S��j �R��dFd!_
��R��;�~@�������J�Y���K��>,\J�f���k�eR�
-2^���̕e\�(�S:���cÉ�׷\@��"X�a+4�T*d<�B�q1xc�^?����A�I'_�-y0��jl#���<ܢY��w�:������ӣeI�/�:��(伛�^)��c�Xo	���z��j�P��U143^�M�ʦ�Dr������섢D�9g��?.����{5�5�⪬�@�lܴ��љ�C���J���wgК���YB#�$�G�o�W"9� t�.{n�AU>�uvH�����%.��:���aۑH!���e�?mP-h��O��L���@-Gu�#����C�*�����:ӷ?b�M����t��P�{�;��~B��M����C�_�j�5��]��L���a=�~�˽_3nhv�S�!d,-�iSx5>��|!k���<H�U��[� !�����S�`�)��(�9a����us"[��K��d�f7bfX�I�cw2�=~�u�p��Esh'�D���Hk��RW�l�) rϻ��U�o��e�.����~�6aU�u(.�0իz�إ�T�!�r���Ӕ�Q�_�)�|�e� �t��S��I�۔r�51�ÿ&�"����Fo6֮	fY�#�>��b޷$�W�~�V��5N�b̹>��Cyp���蛏�Zč� �6Cs=@Ը�}����a|ɻh�Im�)�?�+�{T�;`��Ni���Uk]'�qz�?�1`����� ?�^���k�Du5�>>�k5���Mx�7�/��E�܂W|^M�O���;��4��J����D�ф�6�Cg�G��=w��^��͂q2�,������(1qϋ-��T�R�59_����	3ds����!|�"�Bp���V�
�>�߿�����O_�X�#�pN
��F-!�e�`�|�w^��r$�\,Ւ���r��Zu'�8��J��8�Fh�i dq.�k4�$�N�dğ;rX�2Aɓ�UC���H2n��!�ȥ#���/�欗#���qIp�+��?�\��V�I�nH��O��s�(A��F2m(���Cz�7b�Ǳܴ�:�������Q��\�S�Z���Z��pW`|��������Ð3�J-�>G`��֊��(U��ӊ��a-.��w6����p��5��s��D���ϼ��M������kudI?B����!��R�?�1�Bf�Đ���S�Z\9�C�{��[��ݵ�2=냆���UO���-�_k�F��8h�����%��Up|W��٠���/D�>ba��V'�t9�񢂂Ȗ��gX����*��y&�wה��,��l��|0ii9.e�D��ȸ )�?HX�9���Y����(� _�Y6� h�ӈ��������y���:��0�A��&#���(ަ�+��ɮ�{ɽK��/�N%��t붕��(��k ��9�Ɠ�0�����K�_0.o���6WL��2o��嘀B��Q#<s�.B%q��*C���Iu��J����4�S��6�B��<��gP?��ߖg��B�c�ѡ"<���N��N9�L��V�oU���8^���ƟKټ��r>k�B��{�?��� �q��`k�LD�]ⶊ5�9YNXi�\��R��1*_��=�;�	��i
\m��_��@��Ӏk� :�����xY�1=��[�d�1m��.���Km����a����7��w.�]��K�bQ�7S*��E:_U�,���}D�K������?���('�oTl! ���o��p�7�Ϭx�ې����0�����'�C�Ϛ)Л��i��Br~O��Y��ր��:Yܘ��W-��#���C�'ϔ<� ;MvwMڸ<O��I�uu�-�b�� N��O�:f�&ӭ��6fZvy�'G��,�i��,��vc�U�X2�EvBg_YY#�_U��`�0U���w>m; �o��2��-�]�� �IU��<L���⇿m�:J?��o,�+ X<(`�^�
	�{�J���vqCn�L���,�^6ѷ�zE�!'�TNP���f��͛�� ��2����i���3̳{��!&���&�y�5�x��l_�z�[�����Ǵ������e���1�7S>�b�7D=��'�ڞ\s������o� ���00����|#V~�%ҭ��j�QD9_�����93��o�P���ڮ��B�ȗx�*����ы�+��~ʵ�:*��9�N�hԼ�x��T��̍�r��CH�2-x��3b,��g�,o�a�ˆ�_�:�����[�I-�Q:����v^���}�������f�	�#��:��H�������M�oc���G\�2Պ��b�G��k9��Զ�Dv�qh�n����$��t�3�q��hSS�.�";���ܱA��<"�M*�_���KghSu�ep�TKP��mӡ(�H��n���A^E�bW�Nq_���;�c�XpI�RhL�8����,�=|菅��et�en�,"���uX_N�t�ذh����.}����%"(�YxԼHF�9/3�T����z����OK�*:�Qn`Fe��i��Q%�yդ�����Ȍ�� �>�+���s,T��d^e�k��f^bm3sV��,�No���(uV!���
5��tO�R���T�{Bm�Dц�O��P�Qy�`�_$#B#�7P�J-%R�e`&�~{W�T�,2O��� N=�����|���n[颰i��CąJ��(���W,��jya�<��K1�V���l���vN�����S����z��_#�C���3�g�j��~?حEQ�g�I���(��ރ��ot�\�Ũ��������v�\L��҉/p�%_֒ j���g���������� ����ߠsB �_ۉ.�a1�d�/[�����Ę��)�읆�7M�ͧ3`U��C\���o�)4�L΍>=~��t�ڴ#|&q��D�R�	[���l2�V�ڬ��%ܿZ���O�ɻ[,>��}��ut�������F��i0g�1���}z��ݲ��$�̅Y�j��ZnU�G���cI�0j2�Wh�V��8�s��So����m8vH�$��q���o6�=���BoCR���԰f�S+&trq\
Qފ�H�_3ՠ������SErR���,q�+9E�B
`��;�,''�-�\��u�J~D�	�2,"�����2��э�x_�9���g^V	U���gׄ���x�q�z�h�b�3;�����:N�5�R
�8��SW�G:��/�I K��u�����O��^�.ΰD�]�K����Q˞���C�hf�/ L_�Ly�]�U��C9��\���0�=�����OANyG��S��Y�x6�
���][jm��X�^��;��眬ҧ^I��Z�je]�ϝ͊���n.hCs�>7:�`����g�&
���X� �y��#��L�|�6d�Ҙ�Ŵ2�Ũ��\�0���	삄���U%߈�����E��KU"�2�;v�������!F�C�h�<�4ˎWO�������)��0[?���3�S��?%�!�ҢEs9ƁL�r�qc����;��8yʓ
�R���*�=�SU�1�~�QDG�ON޼ �/�^Bf|C-I��@ktg  c�RQ)��ׂ������b\y`$�z��y迉EM�d���D�$��?=h���(M���U�3�
�<0�������� @�^�'9�d+���q���
CmJ�9_�"�H���k��qX��l�%�{K�6%���A��AUG��y��i�V���@^�$N�)+�;_q��Bh�O���zfm\`���"����@A�Q��B,�7]pQO!��z��$`���V���:��f8�܁���ö����H!(�X����!J�q����K�nT�S�*��'���]O�/�:�YJ�,b��g�����5�6⮢�^*u���ö����/��c�/t�M���Ke�W5�R�a-Rg!���U���o�!ِ��9_�F^������w�m��/l̷f�B�9:)�~`bY\��_�`�I��٭֤k�����M��E�(-���a��b��v<�}��{�;�*p����Y��vD�1�O@)���z�ڵ��i����J��C�DD�0&�6�Ȅ��-���|e.Qk�>"�L�L�6�ըR�0B_tc�@��o.>k"���W���;K�:�}��#/�a
YP����곉wm�%��\���s��*9'�p�QǊ��W�
�����%h¾
�"0k2�͖��Ղ���^i�1�b_N7E��ݓ�H7�z�
�KҘ����qo�.#��x�}�9r�'�fm-[,C���P�R���4Q��Y�	��8�Zw|�<�K���-���M��[-��LZ|7��W��.wP�J��Y"�S��<��6�7vjaTrs_�
'�e� N��GG�G���[u��v�C���i^CɀWq�`����%� b�X4�}B�y�|��� e��g`��]�Pp�����{�pl�F�h ���jB����i�GQ�mvGb���x�=���Z#m�¤Ge���;��@�D.����؞�2!w�S|��׾���%h��Y�v:����beR<�٭l?lCnk3���7ao#N�M�ܡy����{\�\[ko����Nw��O��Q~����9q��&���نR+;-���*L�>�ЯU��-���Q%(\���{�5Q��JT�1O���\�vn�KYL~w�y�!����!K��<#��W�S�TN�HZ��X�5�	4:x����wbN͛�,o��M1%�v_����(�~���2w�rJM�����/��ͨ�R��n������~�9%@T6�emĞ0<��Z�9���Q�TKпf��L6�`s�_��!|�1ћ���HC<�%�pH E����`�ʫMK��me$�cuW�y{Ta�{Ap���F��_�̟̅0E�5o&ө!�Oq+Q��
��n�Aa�����"������>b\lpOԧ��Oz��%����bm�s�
v^�.�h�d�[r�c�v����95j?�b6	%`p�d���:��p ��'x:]o�ő���8�7@���y8���k��p�4k�d���ɶ6*�.�c�c=�,E\��?e�̔_=���n��R����K@�l6.�2j����u�zx7�R��(QQB�����a�@������[+U�w��9����7b����A�h���� }��=���9����M�I?���m�ê���&�3����x9�h'�T�8,niǒ"_��=fkH�]a�SÜ��r˚�k��_�_{�S�ꔾ��ȉ�(m,�k�p��E,��s��`gqX���-�7)��T�,r5��q�Tn��~��27!'Ӷs��p`泀��($��i�'��K��z8[�0����i��a·�Ԗ���]5��F����k����o��s��Fg�=ICJ�,{)VrH(ZBYI!<d��΂�
�l�.��lWr���sUl��on(�P����<-��no:�߭��Z��$�	�)�1�G�u�y٧��� wn�����渻^V?$�L#+z�\-�R8�eg*�7'�"7k�\"&Ĕ�@�[�9|�B>��r�-��ϙx��V-� ���k���4|8��Y�d�Ս���R.js���i����ʾI�����F4�1wHJ
#@�5n�$���Ӕ~9D���	�F����;�1��BN0������G���7�\�SYU�L����$�
��q���������`eI�6�,���x~�6�S����c��'��H��J�NR=A��h�m	Q0�K����%7�r�MR��*�MS���B�h<��ǽ:���	0ٸ��A��5�O���|y8@ߘc�"�����u�he��?	���?[�!��s�Bb�.q>��#&�]�����!�^T�7ߏ��J�@�G��_�bۿ���]-�� ��U�DT���$ls闬S�,��%o��h�(ގ �b�K�ë��p*]C,�_�P��Y����6�Y�z/xw ��9�����7�W�q�U5�bItx�n j�q���R�Y;��T�Dc���f�6Awr`�}�R�SX���]�F0�Kxh%��"�:ܣB����9qi3R�n�~����Jk<�_�ZpB8��}I����1Жu��*�yf ����ɟ��j)��h�o��ot�b{�'X���)*m�NlPl	Y��i��)0�b=�RD��n�H+�(U<H�@p!�����ʛ�]<���X�T�f2rG�._���N?�)BJNȵR��^5�����?�W�D��ϒ�1���wu߰-�G���Ɉk�9J7�z�t0WX�oF:]�Vxה�yp%V��y�u�Y})�\�������� �����2�$��?S��Xn�Y�f��]Tu��w6�L�_�+����|�Y*���3@�� !PI���ި��c�kޚK,�z�G'�X�~�b?���}F�Mequ�* 2�)7�Y5�1��{9��x���~=��)wZ;`�H���+�{������3)��6�fpP�E�����5�6�� cH~������W��ّM����҄8�]e@iXvzA���+��i�E�H�f��r�[&PϽJkI��x������F�����klFW���V������i�W�&�/=m"��>x �Y Pk#�fI8��3��H�p�խb B鸥1%�4 /�����7�}�����Z�kK2xk*��)8��"�[IzŞ�B[C���l��u��X/�?�w$��+X��[*oHtY�K\����D~���b�M��mAx`�8a�I�;�m��pc#ܫ7� v��ÿ��W���ٴ�;D�q��������kf�F��n�-]���6�i�H�.�K��O�NZi�q���fQf�$q��ʂ���k��@o���K��ӐD�S��� M�Ű�s-�e�ϕ@ �����DJ�{;��s}�h�;xNNz/��w�Th��w�g�gD>��j�g�FH3B�m�yV�WU�H�E16�p���%�R�?�4��(r���Y����WT�����(��O�Ġ�V�� L�X������ʑ����jghZ����@EI`
�[�V$�}�,�b}�̳ �,��4[A{բ5t�hcA� U����� ~h��U7��6���;iT
4��J]2)(��"�W�I����Ί�_Rc�1,�.j���3ߩ�]�V�f.��qWh34�Rfሤ�F��9�Lx�9��"�(e���{dg��3�_n"�P��{��!ԴGt�F4�"�l�#3"�^\������;�9��p$�#��g�Tn���R�o`�NT�=��Y��F]���/�>�"��<��ST�OS�Z�eyC�n��ڱU��M%�kj��p�%_(@H��x'xyn�V:S��ȫ�O�)���,1:o�Z{b���{���V��tջt7����d���y�W�Mӽ��c���N���Y!bK�C�\j֣�����n��
��6@������q��\/V�N-�4m��5�^&ӭ�@����`��xu���@�	���L�DZ_}z�3�s�/G�!>�ӻ��#"�y4tb���S{�Δ7�ײ��ٳشP.�2�����۬������6�J�{ee�h�JS����%���� jb�]��A3�M�H>M����4��B,oxm��I��J�>�q�B�AtP���ݦԬ�V�-�n�Q�I�w`}
\�alL�o+&R���v����G��2��m��,����,�:�� Ϝr�a�Z�H�^����l����(ZK�JF����/ALN[[/���Z�~�1��u�\tzϫJ������T0�NR��3`U�v8y��j���d��*�{AL��˴�� �4Ȍ��ھ���]��W1jp����MS&�LͿ�S�F�JS�ݔ��1{��c)�Ѝ�-6�8�a~�Z� D$�&��'�9�N� �Ad�Xܦx P�@�s�5����p_���D~Q�#hx���uZ'�5 Y�62�Ң<��8og}9�o�D�Jff����i�r9`��r2�y��Ӽ�&���;��>��'����b |��L���w���~���%��T+%��|�ʓr�K� #���N��[g�BK���h^dVʔ�"�������kY@�څ�D#]5�h���m,�g�)E�p-��?.�Oٯ��8�P��}���L��Z���8��=�s�̷�'�U��|���3�;���*��Ot-3��t�j�Q���x	���]����I�6k����O��`������J�:�~Xf��v�����P���:|��m�U��B`p�"#�U瑮Y���Ix�"�m��@�Z� 6L_(Q@@k�іA��5����+c��� �W���c�Y>\V~o�`�1B'��K�Y+0/οp�ƭ�(٘��@�alΏd"��
s@�핣���� �C�T�7ak��.VS�OI�����y�Al\	Β���.ݹ.�ӻ���Z��)%/T�v�ph�X[�����.;H��n����j����)�yGfɑ60�gc����������-��˿^=��Q��Y�}N��˛)������6�J�Am��*i,���H���V6�j �vuh�TLC^fx���}{K�C���"ʒ ��%�9���X�yYLSk�!2nM����sʔ�i�ޔ@Z%��W��0����N"4?0�����P�����9g;A2<�P�m���feR�B<��i�¦��Y<�n�iW� m��qѪx���������o�t�3ۃ�}z��-�9
+��r�2�,ퟯ�����T_�b�7}���ނU���5wl+ͭ�)��[@�u�L�|�E�q�\��fքܨ~ը:kL��	nv..���Ua�r�c~A9�O�� ��Pj��l�VԌ]�
��Z4�ìS�H�(k�
�fU&v��T�fnWl�͏#���������{�V�9 ~�LD�X�U���D���8M@UC�F���Ea�!m_�L%WṢΩ�M������)����vm���$��E� ��U�l�0�]Ǵ��1�Q�3���Ww���;���ʞ�Vg���oXT�!.�k�w3U��3� q3��.J>s�3m�G���e>;!��Z�>!�1���z.%��#���mJooyT���e��g}�Dx�7��!2��Y���Y���z���
H�]�� 
��rA�*x�F�et�:Q]5�L%���0&��Ǜ�ҩ��O���;�t&�8���6d���Hgm۟Ɗ���f� g���к�}|&�d/ ꒉ�+ �k�1?���A0�;
�3;� ���J�m�<����6��H��r��G�y<����ޥ�t,ӁV��t�w��K�H��AP>Ԓ��]G��
�x��<S`AD�C8�����Sk�7�?����Uk��+�����dR�`{n����gG���k��%�Y���s�"���r�8���7b�� ��$��b[w�"G^Ӏm���h?j��s�������.?��|ܾd���|�~	 o+m�����8������8Jܻ�z��$�����x���7Y4DZ1Ũ���d��|s��@���Y�?�,u�+�Ł�"zUM��b�"�Ån��~I��t�a�<���ÔH�`[E�/��u!�8���#��E�;��N�'�=;Ӥ��<��tFn�P�m�'�Vh���T�?-
�X��p� �4Q����-v�z��bBxz��<!տȺ�~���)�oy����̨6T����A-o���9�"�Fv��y�=�\K�9Ӓ'����׫�%�U��>�C�	Hu�ө�f#���t0���(1i�UfX�������b����(k�
N����F�|�5��DzT�����q`g����Sv���p��C�8��[��MFbd��&��J����҃ՙ�T����I�i�ıN(J�A��sn��=Y�ђ~(¢��$�|mĄ��ɬ�� 2������u�f��Z"b�����m��Az��}��L�k>�/�Qp Te>Sp�
��YWt;J4ZE;�x�#����T��!�6B��2�h���SK������P Z�nU�Rm'���'�<�|;���iٽ�L�Ë��wQ���n͒*���>��B>�֭��$'9���6ioQ���eb�r��R�៱�l�mhZ�V.Bט��T��'M�UY�J-���ñϙ��1��C�Kt2�{�B�<�� 7�E�뀣]q�c�{���%)�,1��Ѝ�F��M�?t!�"7��/
-'ĵWH��8B
0���q  �4���wcБ�M�����UZ�˿�Oz	�Э =Jk�}V�+��/Ԝ��0�f�[_|)�X'm�x��%�'Hc0�u �^��:3���i��l��p�Ѽ���b������޺?m�l�;B]Ұ���q9��U�U�x�g���~�g|$�i�H���h�U�r�$hϹ�z�+CCG�j�g
�	Țcd�aǆ��ڶ�q�<���.@���ƞ|��PL�|�
w\Gwck[��Ӣ5�1hݳe�&���.X�a)��Ւ.���xb5U��eu��`S"	�`�~�-�#8�����#�_�\
,�03�����%�k��9�^��n {�[�g��[@�Tv.����?�W��� �P���
z.
0E�C�o1�����4�Q7��ai���թP��M�2�T"���⢤��84�A+t���P�n��"�y��d�3(�7?]�~�ؔh�����m����m��_����	<��TR�
3����,v�
��,e�)>+�b7�=�x�,�}� F��vR0�k��	����K]��U����Q<#N�#~��:���&Hyz�o���}h�� �A�yj���4��a��|��ٴ]pM��\1�.��:ro�݅t`0®6+���!����r�x�h��N�!ѹt��Π���+÷�c�SP��c�Gf���'FK�Od�M��~���ra`�H�0?
��� ~�i?W��* h1 �Af��]c"�������;wG�*g b�f�v����#^ܐ�R� ���a�GR�[�o]���h2���C:Xv��_��/��o
�MI�ߙ��E��B4��aε�����e�mS��� :����Q�^��E�����S
��慦f���h@�J�g���؍��$��"��>�lByM��[��/s]oy]���oˁp��g��)ŐE̈��pI���,��#�H�j9���Aϭ�BM�$�,��g��yAT*��� ��#T@����짔w)���:&�w�i�������QQ��qn��O���9D�W�H�����?:���ʴv��#É�^EM�M�
���i�+��ю�+� �$�P�������vڍNi�"�8��?��w�\/����N��[�yͽ�bKS󂜼M֍ �?*2ru��w���6��9��#�NmO�LhƊ��)�ڵ=1pϨv.%�����;O7Q 6bZ�"υ
��4̶���%�񖧟nK�jf~�7��}�nSE���bNl�[sՊ͋Z�S����U�}3x�N�"�R��a��#�0d����	��R���#����l�%�P��9"���q��H�,#=��/�ŵ���m'�ˑ�Ope��7�����S� TB��D���� ����v���KWK��B�=6�H��/���v���m�iƍ�u[����X.��������b�
���f�����%7�>�[m��z���|��/�R�⁲�M*�gb��fjs�p�wn��
W��m�M�{Q滰��>0��Ά9�`����,���gJ��&
J���y7E**��-�@�柅z���c��	�1[:��/��c7J�:R��.��\�
ea���륦)�`n?���R�騨���]h.�{��p��_���C���|�������;v(��_CP�3�q�ṡ�;�px�U/T��tu/sGv���קg���W�}4�|��FX\9��T�%�\A��s��xмd���)�m�]����1�oJ�'*�ۈ���<Ғ���3	͍� T�<�f�F3���#��+���/��h�s�J��h��Rsp�bLO�HW��Z�--`��J�
��h��5�S��;�؁S�G�/��(=�x��-�]��$��Y6XD�����;�c�WǑ�g ����@)��H�M��իHͶ�f1�0�sK5o�+j�2���/8�h���b�h*2�	g�K�f�9�����Pie��r=Rmg>��]���?���|���?���u����J U_�z+3���ym���Ï�%}iر�~ܨ��`/�vٌ̇
l�K�؛=�ԑEW�� �6X�"pmӤ��9D4��l�����i�3����;@�aa\LK߰�U�d���#&��$/-��t���GT��O2@<��zz�����/<�4;����x
��V-0�/�3�XI2@��8~��3e�j�f���P��X�f�<Rf�6-�=�Z�.s�h��ӯ���Z+�r#r���|�Ml�})�iE�&�94y,���S>���)��� l�L(s��d
H,��GOyzX)��h��p�x#"�5ޘ�t�d�o�g��ym���M�d/��=�;����	Tz=_�SZk�UM���Q�yN��q�G�/��B��@vÉJ��Z�_vt�AQ����@�CW�'pכo�m�#�����Q]ߦ��9]��d Ʀ����B�"h��	穾���ů�)@3����ݨs~�D�������Z�|�ʫ�㉻��Mݑ�w�\���i�Q�`��pg�4ITOf/��/�w 5�,)�.��07������6R��v.~�UH&<�b�5F�G���l� A��ڈ�ҳE�i. �U�w�}��w����g������x7����׆�k�A��RU�9�ޟ��0h��a�j������&w�JQx\�O��m�5 f��xx���Db��r"�u4w-��P��6i麰�/.zl0/ygQ���!��d&.���y�r�}[�::��Z��i/���O�w�����=�Ę�jz�O_�������0�w3)�PձY�k�`Z�	]M�|]���Kp�Ⓜ��Q�N	�K��c~�>��R�x�|Ӕfm)7��ϻ����lr�y���7Dujs�+D��vR�S���T�-10�"�ј��R�T{��)W0���E�Md�K���ٓR�Yk��[����Y6�S@g�%L,Wp�7�"���hD��b���N̔ �wyS�˝��1�i���f<3N�'Φ@Ҷ%gr�uuG	"m/��{��fr=u�-�ǿ-�fu֮M`ta��;��%��}Ww�i�:�ԉ5�(��q1�����JZ��gc(�Rs���� 	x�0h�)�7���,���]7�cؓ_7�|e�N�Q�k��T���/E�RK��y,��Tc��n8v�"�b�q�|�m����#��di��p͌9��T U�U��T���"��]<�� �<�X[V��#A7HQ��<-�7*Om1'�G�d@h�%pt�[(g<��@-^Qv<��@�Yx�%�I{S3Ã��&	d؈�v%���D5��A)�R?.�[&���7���9�4x���+��$b�������|#�����&V�}�3���<�b�Lc�}� u]�Bf�:�l�>�ٸ��h?�nyO�O�B�Ӄ�������_0H��3+��|�@��ҳ��Mf�Ȑ�H��4^_�N���Ά�'~q9�4G�����K��(R��n�����r>��[��1�8q�xq�vR1�0Ͷ� 5� ]}"F,�:~Q���K�9}l`[e�=�Gw$��o�Ǽ}����@� P��I���@��4 �\��* ��Z��K��}����a��vb`����gZo�۝��-�ޯ�-�I���NLp��t���[M����U(��8GX���UO�Gp�dc,]�"a4��9������<���Ӯ0؆��΃��~K)�H�p�S��]�B��]����YP��td�q@i�� 2���pF'�bz蘿R6�`���� �'���U�צG�|�),�g���,�&�*�?��(�zeY�#V��W���f�[�ł�6ޢ�i�R��&�=��m�R$G MYzQ��� ��� kt٤�wh������
'e��ek%���q~�1,�J���y��W�K1���h~V�� ��J$����ޕ�<޹�Q�[/W���+��	𤳋z(�fC���4dS�U[nzdo$��\o[�ቩ���x֋���_ `ڛ������`����&Du�'�!l+������5�X�I?Nߝ�|��_���wVD�D�hP�/�JU�C{�F�7�V�v�X�	�J+Ǫɰ�v��������\++��B�`U�BS�&�T�tg����3e�y����S2]��r�;�]���^���!��𥓂Q�2n���ʪ	؝�~��0�L�Lg����LT=13ퟖ�IO��1+�{ ���'�*�zG����6�ݛ{�������S����"�i��hx���Mr��$Q�E����}a��K��	x4�	�4*�UU���%{�)2ҽ�[rr��ۨ���H���&�6�I"��Q�3
0,[���_`8�+d=7�'��$ܾ��y�{09����elH�D*���J�����P��Nn[&�9f_\E2����Uq��ѩ�{G�S{H�Ț��B��)|�7z#`=�װ<�u�Z��1�rp��;P�˄����B��:�z��P�µʛ����-2�;�2�:-���h�j���"��n���G ��.����B=]v�o��ǃ� *d`����Dęߑ �QMO��}h2Ew*!�y�>�����!e���`ќ`�B^���J�X~�!.�A���iM0Kh�4(�)p�;�ܓ���z�����v�9q�g!:A\
JaH �s�ehbV9?�h�0�1嬁
C^��똓�IE�G�=PZ�i-���R�Erq�Շ_*�=m������kp�Z����v�^�w�k~�&j��ψn�!�a8K�8��s��O��	u���"9���o��j�gꍹ:�Y��֗�ߵ��d���D �o0�0d�b�z�veF���ߙ���s�C%i'; �����d'�VnE>S~��ԮQ�ƽ"���֋�J�L�^#HJ��zV��w�l�'"
4h-��t��d
^��m7^kN��f�� }��슾��$�S���*�_�����f�x�a���1V���è|.��+ �'�܄��	�>�ќ�Ӑ-��8px
�Z�ĭP�;�Y}�C(u�i�|&:�V��Q���t-��!�Áۀf⁸p����R�)�3�V�[��\,q~�X]��n�ƻ�+�
5��Ao;��]糸 ��.���P�����|���Ds��f�]c0����;�j �z��g�$|��ݱ�laK�k����I͆���1��l���{A�h.���^R��sm��H��]��D%�:�a3�/�
#0��OV�l��v���� &�co]_�?u�����wUU�+!�d^�B�X��Nԁ;�H2���}f�1���,
�Q��
�7MS�P��Q������W@�pi���b>0�-i&`�9���t�i�/�͂%L@R��Rn�1��g���A�Z��'q-�	@�5	Z�5~��Ũ�m_���4q&Z��U�#��I������w��?��S&%��S�X��}�l�m]�N�s)����in-��9�V���"�}�d��_t)�A���o�;��UD�q����nH	���y����[2:͊�vPD�"f^���gUW�kx<�h)�w�|�M������Qёqv��� f��9�ΐV�D�]y�S���/fs�q�СZ�CH�U�(�!g�6˩�&�ߊ�8ӓ�"Zu���o��TR����
S�}�$?*g��K��j�x���Ԛ���8�ՠ���H��7������'�	�U�|�0�]�|��YP�-OF9�2�Y�*# O� �E��b45��V~a��GEPA�zsc���eI�n�6�eR_��������٤�ycqI�Um�Bw����؜�,yĕ�Alsp��m��zn�~���FU�Y`��=�^@(��.�p6n�t��6�<���.�>k��PX9���t�F��`Z6FQO�<B���OyN��?1_��2�F�J� �~�R=�؆�}�Y��������r�9�/�)�U�N��'�K�y/7�K��̸�E؄m��l��Ѝɠ�j�vyrю����]�k�8OsU��ۨQ{�������Oj��tgp��谝������A-�u?�����X��������
f��H�K-1���~j*�pd����l��,���2���||������8�n��A��5�`�����0��i^��}:����X�4a��HM��g ��c��^-��l	�k�$�F�c+��U	 n�@���p�P�(!�B$q�Zu��Ӏ�Ҩv�T�������4_�)��l6���a-�YIS��n��ɡ��G������S�[�[+iч�q�n�?��֙`�[���-���1��Ak�����Iv÷"�W
�<"�?����bнv6�4�iZ�ն��t�6�#Vq��R7�t<���鎗�:jR��t,�8�l�SAVZ��Ӈ��s�I���0��P!S�&P��X+���jo-Iq�_W��̳�}�Ѩ/m�5/�>����ш�+_���w��֔�ħ�R����([:��+2��G�Xl~v���V�H��ΧZ?˜����I�JB�һX�-�4�����@5[
��(^YC�N�bՐ)Di�.T�
OP'��f�ɇ�Ҡ���:!��V��KT�oI0J��!��u�\(�َ�Z�����"��X#֩���n�Lӄm��đ[�q�w_B�Wz��nW�ýn�D q�p���N�呃�_�yD��� ���n4�g��׊����yD8�����D��kC@܉�(���T��1��-F��P�>v)T�t=���2�]��,��aWWS�����6�����I�� Mr�Ws5����m�j~ �ES��KIO	�|�W������^0H1^0����s�����_�n�vp�����2��U�b)�����$F�]!�Hï+Lk�����8�,���Yn�)�l����c������ "%�C9u����>���ߔ����s����	U��V������:1������M������>o�D�����jֲxY���M���0�\%:Y�X�ۯ1?�P�Z���'_����ݵ�b*�Q��$x�<
f怳�[*Y�����ț����4�n}���E�`�����L�):R�&ȟC	�NNk��>�^���pպ�乆)��5O����k5��`���.%d�L.`i�	�ӚṞҶ����
���J�aA�n�<��ap��Y��e����l$,��/��;m�����W>�~X��6��m9+���_��g0[Q��/sw�F�]��N���؂�-CrCψ'�&ӂ�ZO���1����ND��,�ޤ\����J}Z7+	�U+��7���Yp�a�|6���֬ړ���B��J+�̎�˳��4�H����̳PB���m���WNM�۫:o��)"k9��*m܃W��72O]ظh�L�L$C=�K7�sFw��X��o/s(8�2�֊)Cpn�8�[|�����v����Wv{�<��g�n1]����'n��=lm�{/�t�ç�~�L���Ц ��6Uj>`��p4�[�f�^j�Z]��0劣(�6{O\���	CV��g_x^��Ō�]��O���(���rWl����MU%0`���偟4��.��]����#�Y��I����:��A?#��m��\���ſ�p�cw��\���E�z�n��{W~��˫���"6>N��/�a&/bb�9?��?o�{���-����ќ������=�����2�=H���{7m=k��ȡ��W���K-��w�}�7�E4a^<m
�D�<�3��Br����062��z�P��-x��4��)B"��jW*���1� UŔ��E-䯒�W��q��b�Tӷ,�oB�m��s8)��J��fr6н~�����;���!]����m���A�>&����!;Y=��8#ջ��J)�;���O�d]E�����tE���V��$��x�h�I�i���`.�o�*!�#��ٷ������Ѽx)�.H+��Q������j0�$m	xc��m��i�o]e�Ry����?^�M������q)t#e��6�m��Cz��e��U��`�`n�g�A�"��"bA}g�[CKTSP��(����'P���r��9�Fk�6-fP�����'�8�3��`�&aj��ˎ�e���bȪ#/��9����c䩪�P�.��3W��V��Z��y��M����7�.a�|���{G�[�<%U�;Н'�i���-����. {xd�Q2����c�v-:��3�mp�X�,?�Cûo��j�t���� ��U���Om>/��\w??�
���D����|р�}FJ���],�ze�Y�;4bL �z$��}O������^y�<Y���8��u���:Y���q�ز{���y6h,�v��<�@`(Y��y�i�8�:�JjFXC�;�<:Vhl��]����B3Q]=e�������J�49㦨~��b�@C���{Q@�����R�6ȟ�(��d��hP�P�F��B?�V�wO�a���L���ȡ�F׈������#R�S��z>���J���y�W�Rb�(�᥷��,��W�mg�L�F��3J0�]�͠�	-����:�f/�ư:�!�=A��ų/������&��zc�EN�t�g�qݴY�`q�� ��I��#O��ԡ�,`��w��m]酔ҭ��+QSIƢk���h�wKȠ��M:��3���x�K5z�..�78�1�?��:�RN�S��Й,�4��EDj�|�)1�-�}��hȧ&��~t$�H�QȦ��n��%m�(O�a�~H�gh7%.�)��B��QVɐ�~���2�|�gw8r���R���>Δ�8
u���=p�%���9�ٰ�̣o�3����� E���1`�[)k��F��9s�a9�W��8���nC�ϊ�=q8.�E�Y�T���2����.[�7���!�m�:B���̵,F^��mWF��JD��z]��q8�Rپ� j�e�w �=M;9#��u������(C��4�A�޹K�B���_��{��b�k0��e��tE�O��(V�D|{Ua�~u85k�
�t�E���0�S/ �cq�}����f�[4�E��в�n.��}�ht��]��[�^EK��yj��x�P���A.�/E�r7�ic�9���tJd����f-uJ���C���VJ����g�ΰ��p��ʣ��DRiY7;�i���h�=���0�C���j�X)ǅ�p���} =�3���9�ts{(�G���q�r|����.&�[{�V�թA�`�׮1*����]��۴��a�O�R�ĝ�	'�/w_숤���X�ȭ��Nn�6��/"\͐6� �v-�]�>��5m�@��<6c5�}k�ńm;4&+əo���x^�[�lђ�z����HI8(z�L�@o~��
Ś����U�?��Z�y��ʗ�m���5H�ߣ����r�i"�yy�.яx��6	zCW�6[�����ra6�7�:��uM�<���v7��ٳ1\��*0Üݶ$�_\��C& ��µ�J�%��gG���C^���H�(�/�����!t�q-tm�ǃ���H$�+4߫ �aqМC⍇���ǘϮ˵x��E|C�)<�;�A��v�]�xEn��e�t���甦q�,��|��-�)�\�N_^q�s2&.���iaX��d�a�$ .����D7�謗�X_����Z��Tz�4��\��Ҳ���/(ݲ:�����)w�S������+���%�Z�+��{J��]�n��Zn `Oں[^F\�P傀�L{>�{�D�Os('�^ܯ�V|r��Dy���t'f�"��RYO�O:\�.b�$#�N⁆l�d�w�����!�EP�`��k����0b�^e�V��a�|,OD�m�CL�|yV�_�/�Z�Kw��ݶ�,ď�ۍA��|z�����>`���fW��]��Xw���I)(9���\��

	���a�U�n��T���١2H���&bl�pSE��u�n1�ev7-X���(��P��Fz��k�d�	��^�8�O�?�2�4T"�ͽ�}g�m��O�RZ.��ǻ�@j%����L�Ѽ��-]zЫ�QT�A�/��rw��l�6�[�R�5�����O�����g�m��{�l�\�Nr`��;����9ȟʅc�YF6\y��Gɑ���F�p��6:0���F�a���C,�8��I׾���w��㷣���)]��V#{A����n3��&�s趃�`��~�J�p\�:?-�8c-��X��5��\��Ә�D�B(�|iѫ\��#%6R�2Hy?^�(8�3�/���{�t����i��X�g�SN;d����_�����-i 1��#�(QQ��}-:S�œ�^���w�tFIٯ�O��
B�u�[I<:F�g�����v�������F�q�q�"L$EC��2ϸ�`���/�`�/�f'��~y�SG*��g��0�]wԏ  ����]�b�0���:�f���q`�%�f�d�&�d�|w��͸��khb�R���0*�3T���:���upi���|@�W!��Ze�o r�	��./&E��2I{ ����;f���c�,�nS�7���߹�<?,)�-4p�@�4��7C�ٷ��%���_<�m�p�������DZ]���r��q,F��Μ���4V��~�N����G��*~���p&�59o�[`���nu���tv$�w�HV_:Ѓ�.j�u��2Su�$W��%l�~��S��_�!J@�m�n4�%�` [���Wc���P�G5Ç���^/���� ���d�kB#�ʟ��H�*�ʁ�5����Z��WɡKOkh	�L\C+��5;���\�Q�:T�uy��KJ&��U9C�@�<� ��f�d$������)@��/���!�W�`�b�g
����z>� �P�R�r�`��`"3x���� ��'�H��T�Vc[�r���`��<n�ݦu�wڝ.q�Ji�kN��_(�0/��X��q�K >�y�K�F^�]a)Ʉh#�
2k�0[��M�ɭ��ԋ����Äb�2�y�rڦ��0��l�I�p��=� ��撕��kRi���w��7ٖ˝������Gj�p���m4f�� ���ܜ��r�j� 	�v��؇>�F8hel�5������=:��+N�@e�R$j��؍z�I��}�0�ݍn���y����S�Bn�}qN(�sDj(��0(��Jw�j�Cu�r� �z'��TZg��g+r&X�t�h��!䣧�O�����|���/�<91*�%��`��JWv��G/E����t����~�.����ȉB�ఞ��w����g�r�F��[􃼬vz/�ΘH�]�3�����Y��͟�JP��������İ���rWa@��oXB�c9����;/Z��d� e��'ݯ��-�Xnn���� ���4V��~�������JxĎ`e���+˔G\���
�hQM��Gޙ��n��v ��ڰ�R�nKV��v� K9��@�A����L\�&���6��MPI)6��c�v������]�{��f�Ht�F�n8ϒ@������W�H��sm�]�4�J;9�d�����P�T�S��j���R�{=���e��
�j���z΄�����x��ϴX�TA9�iˊl5�Gzd=	E���L�2�,�v��u�eWC�&Hc�Z��z�HR��㯫��܂�<�.j��A[!(�{یʹO�c��C����J��|]q淝��lr"x7��?l���8b��$S�V,�'.(#�E*-f/"��9�TW���~��!�w@��((�&1þݓϡM�acSD"��x�~�&�9�D��\!��SR2E����@L�N��Z[ ����K��D�@�<�RV�a��I������9�)�ʏ�\��P(L3��&��,��s��"!����vW�jE�K��jR^wx��������K"������]yX���mI����%L(��-��9��C�;qCc�o��)��0i�$RSJ|v7m�ط��n�n�`�$�N�R"!˰[ͣ�X�ֱ�k-ݏ������#�Ǽ������!����@���A�r_w�����>(%hI�������+N��*�d��J�����A����v��m������u�/�<Sg�'�a|,�p>����@��f䬉>�^,�0;�T��bQɑ�S���JGCW6�k��}��@Լ�C��n� ��7������x�<��d���I�V� �)����DB������XC�F-AW��g�������A�D|iT�h:H� M.���_�7#��HN��Zj�k�@�9|e�Q8r�HN�����	K���i,'���V�C�u�ug��@x��%S�B��_+v5&�=&L4�<�e��乑���E��{ڋ7u����A�@����'�ހy�F��Au�|��V�&��(ty�7\�5�8ZO��j�� o9f(����@�PM���'�2��@���փ˚s��]�chɛ�֨��"��>�K�d�Z����nP>g����W��!�q:��e��Lw��[���e��i�`����֣o��{��F��ې�L�SU6������^�e�P�g�'����ӎ��}^���l�:m �5�k�(�����<�A�����/���I��|�g��TB�x��.�"}���[Q���n�wa�0ÿ@��T<fߌ����K�8F�N �5��$X/��r"��Д@=���#���ͩ���Ē��N8��o�s~�
l���0vD��XT�ߋ�ĉ�?�-Hh����*{�:�+�wJ"�7���B�vwf�-V����^��vY)�P��~�]�
��C���{J�
��#�"��Y��:�*eO����[u��c��������ߙTK�V��F�~⨦�a�SdE���3�뻉P�E�븸�ic�_��*�N��@�U2��)�l@����w����FZ�h��W�&�:�u�9�fB�d� �2�h�o|(�.��M#�Y�P�a|�<�����ٟ���2),��P��̞�'Ʌ`(�Á]͌7�?��� ��� U�_*�A>����3�!h9��(Z�Ѡ%	�����xփB��<2�/��s>A{$��sb���#*:�)�o�b��s�[���;>�ۈ���P��ܕ�m:!4|4gS�p���_���7��>u,ta�:͉�l]�K���ۓ�N9�(��r �8��Ń½V_��і�ޅ%/Ы��/�{c��c�̖�I�ws�������*�������M�p���xL&tZ�fv��W�vڪJWu��{�ϱ�K�}�[�hEu�y�b@��	c�'R�:�uN:�Ò��ԣ�y�/(�Cj��L�so�/�ׇ02ޞ������ �S봗�m�������&u�p?�DU1�G���L�����!bH�F&Rt����a�l0CP'��S�ZD���<c��Zw4u�6��J��H�&���'-�Ds*�1�A]�?Y��Ye��F��D��{9���t%��G�a9�sh�c&t��WP<��q��~W�<�����ӽb�ڃ�h�}^J�������d�DV�8��S&�<��8p���V/���8�!����_���Z(0��YL��1�5d��-c>hcWü$�iB1s���6`=��众J�&Gح�ɑ�đ�q]�{M2~M� 0�x>����c}���!Ώ�r����r�iU�!d`FA��Օ��|����%�Svϋ0��R	�]&���We4��9�xfS:�2)-�s�"�bh8��^($��nO71z��+����]��:��/W?�	� �dY5d֔���P�Z�)%�]x���O@��K�	+zI���$��h֒Rr��S�,�hi�W.�7�\���&��޶(�����Ɖ6�QÚ��ȃY,�P��st�/d��t��!`܄����ט���C?/k)B���ǎ�Rj�x����C�y�J���ğ�u�݊���;Y���[��j��H�!��AҾ���S͓�a��P*2��`Y�M�k�eT���:L�oX��5r�3��ё��5㼲PQ�ى��91��51�e>����B��ra7Ҵ��H���ϧ�݌���fr�m�ծ��duJ�<��b@t7�Ü�6��]dd\/[�kn�'_�NvwQv�"��7��Ղ.�
z�w�`(�����#���>R;�	ԥD���CH֐��&G��Y<�LH^���MO;���ղv��آå�)��n7|�~.,W�J*VN��ֆ]����&��-�Xw�╧f/9�EJ�~�h�«����IŒ2ܺ�!�y��L�9��W�f(�D�4�u�j(�3�G�x��+	Q��w	�W����׼�ܐz���9�o�A{LƫK�,�hO*��/�����//��A�����e'p�8H�Z�
p���I�8v.$0eO۞P����mN�ؤPŵ��4PYb�z�u������W�!��kTu�,�����Qx/��P2"���(��(��O�zj��9J|��:3��uECҳ�D�g@�ɚ@������u��I��|
�������meW�|�`7 ������Տ+���~��Zu_�ON��"�X�P��d���]�I��,��tC�	6Wj�(���dg ў��\��f��i�w�j�J>�G\ѩZ[WH���vsc�C $i�!CN�ZQ��|��O�ɂ�/Ջ�@�����he5v��f��5��ܭJ���|����o��q��S�y�:p6�d"��V��cb��x��ɮ-ŷf7�^��_�(�;���C��^T����T"��>�k�5�����6�쪋?�>��1��a!�5����s�¡X�-N����>��{9
Yo��a9��i ��Ō�u��.w�\�hmMnC/F&W�y��5۳�F9��Ln�	[`=I��=5��D�fd�;�P}��,����N;�1���],qW������`T�������([Qw����~�¯�+4�
G�;���=� bʂf�LK��%@[��#>o&G�I��^~��T�PC��@�Z)֝����k|Ȓ�Lg���:ӈ�6<��N��۽�J�6��e�T���n*�7;&�R�#&�m�-(K�l ;?Ь�Q�F�G�$��>��:+����G��E���x�!�=�6��O�/���Y��L�-�L��d���g��&�߆B��Z/���l7���8�հ�������]a�nl0����>L5w��k��.v�}V�?��j���6�Gpu��e���GG=ڬ� ��nc��%d3��8��ea�L�:&���=�lU�{�?�E1�1��9���
���v�� ���3.�#��}V�̓�nw9�^���E�.�����4��z,��h5��n�d�o�����F���H�6?)3�(wK#���:������v�h�l�q�[�E@";���3ئw	��7S�/������|.�Ò\�W�/"9�A�!�=��W�5ǃ,2J����U	��D�l�U�o��+�N9|nvo����t��/�ë��v�Ue����*�(t�e��\z��`����l��G)ȰAϰ�erK:�[�օ	���8L!� ;.�
]��\^�yu���X?�����A�`�Me(��^�o�7|���%M-mfV�� �@z�������=r�>2$��m�JJ����_���&�>{��А�
֕���$Y�U�A��e?��2����3�+��qSS�\�tMV]���q����v�h�$� p[��3 �:�9э+��;���j�{Ss�).�Ə�\�$bђ*,O6�w�j?� )��w��@*�����>I�5t�Տ�0.N���&i�� ��o�~�z��^ ���<z�'�)h���|����]���1��-y��P�U������#�N��rR�I��D���2[���*�+���=�j�e�蟤@�ۮ��3xL�p�6`�p��w�8`֫�z�'*P�� =u�l:v�JkuV@!�ؕZ�q���٪�3N���6�N�\��v��c�&��k���{9Z ��q�l[ݯ�ele{\y*g������~���E�\U�"`���Y:m��l����*L�{T=pc9��:e�d�vS��t�)Q��Y��^�ٳ�N*'�v\�dr�����WV���� ;�7k��*�$�P�'�>m�v�T���N�Ke��&@�v��� [�k�p���zWż��zQ��j�n�؝�*�l=j	&,{;���b�P����<{6�b͇�3�w�%7`���}��d�>�9 f��*W�ߜ�)�Sh����aG�xf_Ba&�Ĺ�=�X���h>"��{,V;�iIW�1��$C�������KsL&��Y���9�w��<�!�7\{��4H�t�w�j?Uϑ�t����d(gC�}Q)̱�}���R�T�<���5���DFk�q�����Y�!�A���:i�v�C9�oM���6��A+�΁I�f�;櫲��xc�&e�z�|�c��	z�/�6W�z��?v=gGX�m�l��o<��eQ.R8�$��z�J�v�Y-��Rǐ(�w�:o�m�x�o^�ʠI�&��x�u�����\r���S0��G(��C`��_��kr���H�<�в6�z�R�QBA�$H9�Y����}/^�wbVbD�	\5@f/�����y���BL\^����28'��߂�W����$t��k�z C�er��v�˞r<��l)V-�fg�u��9���%������n��0�?����3߾�$���AqQ*]l��#t̕��D���������}�� �X�8{+3����b]>�\]{2�۔n��܉@�g;22}��2��Rn~�*��A_-vD���E˧�g�~~�vg;����n���H����E��:�����Q�1�m H_��yr�c�I���-]�3�q窒o2����'�X���`,]�6�c=��̷�D\��^ ���,��P�`7��Wa��&�k(m���`L��izE��~ٔ�M(�QȂ��%�/eCCv(��T����ł{9�Ȳ���j��Z���H��О��.���D�<��1�v��*�ޏj$�Z�Nu�6l�h֔�x�O5?�W/�`��K������[��c���R�^��|R����M�x����P1��ϙi�z��]�@7�bg��4�s�Hq߼J[Ҩ:�j���ƝRͷ�S�v����E��C���} F"�@��8'���F���R%鴎hʃj��;�n23�&m��sA�gП@C��P5�\�dg�S-�!�H�w����.�E�$H�O���G;_�q�W��t���w�쏰����H��hP�P�U)���ޛ�2�|���w5�x����n��GD����C0(���e���mD�ɕ"�ȍ!��r��i¯�D�?��X�H�Rp�.���$@��z}���E�h�r�@�l!�4���*�d�MN��+�G�;��� �O�wq���R��-�4VZΡͰ�����:�V���ѝ5`�y�p�I���I� ����=��4���y��U	�X ����_ԱN~�)�t��w�/:#Yk��m�1A�ИD�GL�y"0���hi.'�9���x��I�tc�Oj&l���U1�)Hb`\;:t	bJ�A-e�����8��Ϛla�����x�k̄Ai��h>�z>�|�y�6�W�k7 ��	�3X���M<�4{�*�u��1�X{�q\�����.�hF������i�p��p��M([�<��>v']��Z�Q�����S�h���0��y)H8qN��o�,�^�g~q��:,��lp�DqW�{�?������n�� X�	@q����3ylP�x�6��;m�Σ��2k$%ӷ|�w��tx'��.I���5A;��Q>ᖝ#4}G̵Ј�$N���+n	쨝ڱ��Sg
�wAH��|~��y:��8�,���4��7�u�_�j���m��r�Q�D9늲�Z��&����DR�l�k�����R�]�IΒc�VC�mLg4��z�ȍ����K�i�Xm?d)�;�<�����ss�q*/13
ݳ=]Ef����13�}֯���+����4�@E5��.�D��6>:D�}�H�D��4?Ҿ�u(;"��o�՝ /H
�Y�QR��9�~Q/�Ͳ�I��� ����Ŗ�a�\��E�8)e��Ɇ�A�@ٖ'���V�PHg��B�/���*���F�l^�,�`5��:�0�R!��V�{��oϩ���<�dT��(n;�i�u��w@a��� �ŧk�2W���?�ŧ7<[I���h����?P�+�y漸�l�U�^��q^�#@q"&E�(�����D�2VcD�G��GxY��ؐ��uDɃ��T�G�:�Uz&(���Ӧl�;wh=hG�Uu�{|~����P�qJ�_��O�wdlv�4;ɥ7nb
)^�)�CC<8|4�g�������	����o6˾���P�ŏ�"0��K7�l�p�G�ɤJ�<cN�i���J�oE�-��
��;���֤�z�zj�n�x"�գt�BdY���v-Gv�[���#zT�s���w{�h���6<x=��\���|�o��K��
?�{��Q�����Y������zR����>r8�̾�6��q���'�=��S�@��D�� �U+�O��^�s#�b�A.#�Ll��$���O��i^�Y�NW�x� r��UĒ[Ӕ�a�R`�M�XB�v�Uf��	B�6��$E�6���^�K��?8dx���_����ٌ.���P��:菾R�����d�l2 W�� ��)���GD��v|}Ս����OTY�I0��k�ڮ�.�w� �nb�c�����̌���dYߕO���GVD%e��+D�7�ݢ�����Y)TNE,����W���~�a�;M�I&R7Yk�h�����s�2����7f��Mh�B��&�!Q=� 5��8���ԾVGp+B���V��.y.p�e=3�Y�I7W����(�Qk&�1������->P��T�S�-m�������2� ��"��k�԰��2�)�������d�Ln�ۙ�dakY��2��*�MԖ�J�^�:���n�O.��Ƞ�^��ʮn_��%�)���� ��!��؁>�,�#��B��>�y�*��e!�馡~�0��	�+%p��+���p.W���$�.M�[�ߟ���t�k�&.��-���>��/0|2�m~
3���r0
�>����G�Pj�97��L�Y^.���-��v�'k̒�ƞ�����R�,�ܣ(�w"'�[]�:j�N �bre]�J���a���^��]о&��A�,����������}�~�/��1}(�|�K��ț[�Sq���n)���s��.�e�,�t����n|��D�"��+@�K�71P�xf	04�8�2��Ɨ!���Z��!*��1�U�;tsوw�.�Nh�����}�ٓl������쁵d��'yL~�?����a7���@G�H^L�Fm����>z�h�*��Q�����1*V)5�6��[�._G*��D¸L(�<�`)��R`|'���g]�xU��B��:ؕ�Z4�ҫ}�K]=Q�&�Đ����Y�[<�VU�8�S�#7,=q/C�O.�ݺJ*����Dv%�	=�g���~�IC߾)?�WD�F�l�����H"�VC�ɶ̣���X9%�=Dh�2U� 13��!U�2h?߀M�D���S���Ҥ��]Ԇj�6hk�ӭnӪi�+nH�����P�r��c/WH�Pe2`j&d��2��ٞL�I����w�B�v�G^
�X�j_~��-+�!��+��aw�ltl���Ah�	��K�3@��w�������[Ze��h���N����[́3��]V�$���C�{��d�2�0�!��?�GA^�Ks���;=��]QL��H��<E*	�����]o44ŀ�ۣ��A2$�+Kw������B���|�=ww�O�)��К�q���XF��)��v2���V��*1��m:=��@3,�&�c!�r�E�'_Ȏ�ng���gG���*�'o�)ݖ?'�#0�P��F�'Sކ/�ӸV��#�IA0q�b�u���0��3��G�&a��4�7�X�Q�.ZDbH{�~��(��*X~ mv0	��t�'5�1�F�/���F1�:"0L��Ts�N����n�&8 Y�$b�!���m$� �� M[n����5)T���tu�Y)�ЯHEd�	5��Jp���N�\E�ӹM.�9N��Eߣ{M���*���*V����I�v���8�ڲA�(�5r����|�iK��{��<fF�H��)tǱb��8���_H'�1����t+�;hla~�.�A����f|oas[��#Ke�ud��]�EP��>-�)����Q�g�q�IםbXO/]���s�/Ox�Fv��C!����d[&��<��uS�x�w��17l2�?t�nm,S�Y3�[���J?-z��{�P}[NQ���	/K��^%6h+!��_�2�N�N�U_cٟ���mm��Cɞђ	��ݳ&�Djci��݌pK��ɒg�M��d��_%�&�i�,O"(=D���ᒤL^#H�L��mcOk�w{��I���F�N�\a�M�#��To2#+�0�����'pj[�6���(�7�7�,6��c�n���m:���x�y�	4u��������	;d����\�w��Ҧ�׋��홽٧���?����ȋWCY��d53���y���u�*�U�1+d�?J��(��b�?E8����"��#>s������vJRI�l�[4�RI��G� F��$M���wu�og"pBs� �H>wN�\f����$�?��}�۬�C�o�~y�nWnkI����7��0kb�� ���ƙQ�O���f��"z�gNnoE6X-��SGAT����11���0;`�0����낹�!���$���8H��o�9�NĚ�����~%j=�������wZ$�SD���Զ1�R#0m���]J��N|�0V�%D��|֚�w��L���o}�g�	>c���g��mr�V�k�6�O����!;�>��t{�Fk�x$���|���BgCm$�4�I%e^�		{vl�]���9G�IA�����!��$ۅ�+/���L[�#�؈�� K�ɥ)��5N��G웗�ԃ��̗~��-j[�9���m;��BVB�%l|w���G6�r��.Z��9����@��\�{�0���@�����ǘ������r����.�;`�ˈ��gH��yƅҖ���9v����ue��i�[��hǾ^>�2����h��+p���E$-��n�����P�A],�K��1�bu{J���T씶A�$�4Rdײ�-cɍV;V'_#W���v)NXkY*��?	�;=]�c�&�塘nuh-�-�8���#�&qɺ��Z�^�{(�hƪI6���%�vqm*Ɏ���\�`��#�T\uJ��n�%�|݋!p�)Q��<f�u�Zs�(�n���Kْ��C�n#/�6���EG4���Ȯ*M��g�@y���x��)�d�
8��C��1~E��W�rv2h+�,�IA���/� T�	'5.�C瀐h�t�~�M��#fx�">�Ivϟ���GոŢ��a$��2�X�I����}�M,�3�9�?N��(l= ?��b�X&��͝�e'4�/N�&~&2!��ݫ�l7a�ً�z�,C��VAo|�#�]{�τ�p���K;D�RMh�KR��v�'��R����	H�����0��g�"�~gb�=:��9��_��+k 43:�7}Y�:���ƕ^x*r:m��m�椪��&+�p�2�hV�﹭S��dt+���TF����������g�w>S8ģ��v�d�ۿ
���p��:��{9����MH���c�*���͞���4"P�`�͟:��m�L�r#�`�n�\5i'>���R�&l%�Nٷ���M;�6�]U�cg(g�´��g/���4�u�ϐ��J�ړSL-�`�3���4sN4�J��=y[Ƣ~K�Ҹ�[h�;�)~w^������G���n��m��2����grm1
��XBmoT��pkNZ���kg���O�����Z[bG_����_�@����j^���9/@ն��u�V׃�o�̬11��d}W
�i߭
5S�� ��-�����(/���j�B���h*r3�a��4ъ�b3��Q=��¥�l��[��[����HX�����V��	h��$My�E������J�U+��m5�0+Z&)��¬�;�9H-�_��d�hdk��.S^ea�D�>G�p*l������VJdM`e!�wJ���B�M�F[x��Q���;{��s @����ˬ�Z˳�pn0C�T������k�h�������<�!���_?|�_-�P6{��2m���E|�5�q�p�)q��7�N�(�ɺ��o���&9U��
�ƣS��2���
�&=���دȵa����.�EĄ#LG���������1��Ka�ؙ�4����%z�.�ۣ�aP��L�{?l͛�^�d7¬]�����W��X�_՞k%�u~]�h�/��D��l����<�¾��e�V�Q&�v������&��}��t�JZ/1����l�S����_SH��O�C'*��HA#��=N,f�B:cǩ��'d8�� u%C��� ��e��L2G�`����f>�iCD�ڌ�%n���a<���[��jT=K`�8|G*Z�ϯ|���������Dl�+��Lj�(p����V�G�6'�����8��MI �V�рKB�p9"zc�sDl��U���p�u|��Z��I=�oL������(#"xr�B���������P(�;�H��6/6Hp��_�]�����.ׄuA�Qw�4�;�M�Cp�>��A�8?'n�k���ܳ,G�k�%O�j[�����Te�<�}1�Ƶmۜ��ذ	��*�9����(LA��W$~(�)���iIx*�MZ	��ERF=��|3��%7�g�b�}���nygR�2���:�C��+.�qT����4L8Y�������c��� Wc77�J�AO/�v^l܉Z#[*x���:nV����7ϥ��7��II�r�0n,�s���������Y����Zq7��_���EcWc��f�ep���;�|�vu�ͫ0S� �V����6�h�FRSť@s6)��k���s��W�	�QdJ3&���:�������<yu�ח�����F��:��#���b���D�'��˚�@Al�0L`%Ǯ����[k����g5��E#x� 4���P�BZW�����1P���b�{@dV	�N���Dxѓ�۔�+�R�1�2C�`/�"e#��Ʊ;/����N&��
�<�&[2t\���I��U������%�}����Bih���=`��G��e9y� �2;kvUC:g:��<"0
��dT���U�
8�L�	5&�$|�p�MY�OGd�E`�	nr�ﶫz�8ȝ��W���ռT������땃����_g���ؠG�1��B[� ���{~��b��/�g��پ���w��m�c�+�ENČe+k ��ȏ���/��n�;�4��.z���+CqWV`�[C��V;�ߠq���L���~�����' Vv���-)o۽9��s�r7��M�q���R��5�|T�;NC�bN׼�fSv�n�j_�eC�J�1���
P��XÊu�s/�[��J	u{",;���@����)��X��^SF5�����(�>��4~7:`���6�	�J����Dz�9�����+D㸒`w�D �/͚�T�]��[��.�)ʌ�<�:,�h�z0�K��W�m	I�X+@���˧!E/1����C;��FA2�s��1�MVE�8(��1~���O����j�F��ɪ]��h�Q���
��Z��Ձ0���z�R�g��8���^��N2�Ҵ��9�W�ei���et۶Vu&'�
0��=��~57����	�'(c��^�Z�._���!L�_"i���2��~Mҏa����H�EcY����<aRT����H���b����/���?ly��������/�k���nD��)�"����K{h��E�O���v���{qC5� IQ�f�裣�ψ���HƗۧ�VF�a��@e6Ѧ7�i��*�0%����/]��x1��R��r�;����t}��B�j���n�0����;�f��{"~��W�2�`��q��b�^���S�i�ق ���Y����O���0O)�N��dӏ6#E�"�;�Zb[P��g$��6`%:����_���ӽ�����'��0�a���L�r������l��� dN�q]:��v�h_�UA��2B�k�4�y�[m�ܩەo���('R��.�L>��ߔ�;Lv���bI��8�	+d�����A��C�`D�1��KQg31a�g��h�������z���N5��>ҏ@g��G(��C��r�0�F�
�,,����|�?�&NHre~ru�Sn�2�4�9��Ѳ��� 1�tĖ��d'��M�T8�0h3�A��U����:,tքV�r�c��Y�<h����@w!7q�'>���j@[y�f�i��I+C'/��o������d�g
3UM����[�r6�1(�q�/�v�ּUmCG�(�2��Q�.M(�f���]j�b��B�!Wf����	���iWz�w���=.�	Iװ��F/=�5%dgIB�2��v���V{9+3t��Y�_Tm����?�p~+,�Bc<�_?'�]��))b/N~���U���4���+�Y�À�FmK��h�KJ0�e<+���������')�e �ǫlc"�2��K���j�Y��ʋ�iכ���[O��]��~���:PY��X���bRz�Z�I�8��g[�>�f����#��8B
�q��6T��NFGo�^׽����O��^�ĩ�0C�� �r�SU�U���j7J}8	0�}�-�S���m�C�:<]&�Tk��9%�E��<BPӑ���S���e[3���2�64������ �`�в��P ~�ܔ�;�-ϑx|C ����X����D��d:�H4�E�|��K��<8�IJ��^l_�.>� ԥ-�!k��<D�,����ޯ��&�[���]��T[Q��4#�6�����"F�f^=�.�q2�������e5q_��[2=��=�0_�ڑ��#��_�ts��e��^?�N�Y7yp��"D�1rd2b��]R�E�u��w�n��Y���}��},uu�x����z��ؒ�l�;\���'��ݧ�P �#4�"�좰P���ڊ����FC�r��=o����y��-Mr/xq��ӻ��=Y��%�䙋�d���6�� �̨צ� ��}u���>�y��P�ھ,��'��W2��,�vFg���*}��n	��@�v4�\�8������$��w�K�RXG��$�������Y�_�"�� }"�  �pY��*��dS�g&��6p��2�֢"��,��>��@��r[d|�w��mG�j�^N&�_c���Y�HCh�Ok���2P1{ty��?��Jm���t��
4	�mݰ�>4Q4�i�~�э�!2�Z�����w��Β�T��a�6���I���wz5�.O��&71�Y�w��Ɉ=�j2UIK�Y�����4VZK�����8����s5'i)�����0���8,�q"R�����,�;?�y��V[A9>�����zo�q�ߤ��(��
���=�B:U7���ȟ�E^
��,r�^G�B�+֗3���J�E��ਕ����8�2�:�$��??�i�G�K��?�����37APht�,i�n�S]?ނ׵�ĕ�s����_��U�gP�3ק �4�X�4�a;�8?��^�$
m+�N��X�Ar|��_�J0H����;N�l�p?�~���%����B��1�`"�&���u��H�R�ϓC0=�~7���>NM�49%VhD�S\�u+�}��Ho�����zZ!�ˊ�wR�4i�.�>ҝf�v9u(���~.��K�G�����6Q/4&��Ɂ���0b��/7��V["c��Jz�?q\�^XC���n�N�g�q���I��go�>�;n�odB��ҫVM�U�1lhݹBH��x�)��b"|��G����Q�ȵ�U�;��U{� V�z�!F=��p���\�Bc<�43�o�{�|�Ru���=�y��QDI�y`u���cY\lC���~�a~� ���NVNh���jw*\b��N�Q���9�xC�&SJE��7?u`�,`
�o,��;�������ƽ�=�B�6w�Q�u�h+3�O�L�J��"��P���+ޅ"��:�Lj����/r�H��&���m�ly�id�W�&^�K�ݣC@���W	+yy����>���~���fS��������)$D������=:�%�9\�w8�>P<yQ���-���M���:ga��͠-�C��g��Gw�8L aMz󿵢7`�.m����#� dx��:�N���C�<M���⋙����<�&�����C"� hۭ�l�:�G!��$Z ��+��
j�����}M~�L����OqM`4���G��՘���2�(`?NQ�V�+�E'��6�gB�흏����*@��'("�_�?߻���pÑ���E�G!r	}�[0\�뮷'T����4Y�'��4�%Y����t���Vm���l���.4�y*�s�uƃ<��m��$��Kl��_��w2Gv�]y�ܹTraq�����!e�q��`��}@(g7����(��=x�W�{���4q�\H���Z+3��q���5΄��f�)?�����7��
�����-�ZS��&���u�c�郐$~�� 5��=�nyt}�z�[:�j^!��Ԝ!pt�?�?��0��zf!?"��>!������?�߅/�T&t�bwNa�e�F���c[F�PM�8�t�XJ�]]D�T�\>ߓV��sS����y�̀��`�DQ=�b��K⠅T�N��[̲��y����nv�Z�$v`�V�Ie�bS��y+H�2����;XhDܭ�]�h~y+��8^������c�	�h<��8x<m� Y�(�灤��5$�&���O��#���
e���RۡU=��e12w��%�U�P.g'5��o"��;��n"	�����=T��waG��9$�/	'9x��!Y*ӎަg;���"V��� M����hGC�ǈΣ(���h�߾+b�T\�;�J��"��������P=�1ƱX,+(��{̩�>�v?�_�I�7̑3���чwh����§���wp����Ӡ���+hqk���)B#��C����2e��Ź73�<\54��j��i�%�����r���xX3��{�j�X.����7��@��PEuȹ �R�`����'��� �	�(t>�ӮQ�Ծ{>_d_Q��q�ok�6d}�������E�BN^�`����{D'�[���	ƍ=0]�C�؈��� )P������7ĔO��{���ZY��>�P�=����lR�_����Scԝ��:�t*4a����P���Z������n�h{�/�Gw��N���I�>��И�3{�`V2̔��xJ��|Kv��P[.���oc�a��ݹJ)�FĖ>��>�I���ܧ�rkM�E��}�� ��:�s��%���ʒ�@�A �(m��3V'�JIDMd��W%�~~g �o�����Mr+ Q���gW���j�!=x�E�/�/�����]bZ[R��L�A�`��N29)N0��_!l��$V[����4M�z�^x�r�\[��\S+�n�^ �f��
9�f_C!T}>[�[�p�1��E�F�)���U��1���ep������Vr�1��Q�:�Q�[���N�cb=��ʞ�FI�����	��
E�*��46��^
�&�l[F�iN�D�X�:2jPR�DOP3��Ӷ��J�<��gh�tp��;J�����!��7�`Fm,
zYv�m����@B'�Е�3,Eq��a�.���;��=K��K.[Q���Pț>�Xḋ�E{��`��z��nw�\}�->�)���??��k�jW�M&,�����X�N[?���iL�h{�T��e�|K���ɒ����-(+��j�D�p�/ 6b&���23�IR��~g}O��r%�H��XC]��)>�`�(uu�ɭ��a���3� qr���q,b��z�
�\�==huEy�Yp�x?����ɬ��]�q��%t����!j�ǉ��w ީ�΍��5�z��Jo�Z5�����Nc���9a�`hPg
M
;��q��r��w}N��hmZ|��۽K`3�6d"��i$�����7���D>��ZlM��#�}F�쭙j�ӓ�rk�oZi�����e��{	5�r4v��zVO�����9��a��q-INL%�S�ix֍��YΙ�}f=���fQØZ�.�"D�{-'3��&Sfsn�[��� �7Y����켛j�!���U�-�{�!_�?�C������4�d& ��yH`���������TҾȎs�d���V�IӯH]3��(H��)�u�KA�{�#S4=��C����)�zǔJ�P��,Qa�Ж��L-�f�
�t���{,��^��c9J�'�A�!���:V��2R����*W_pq�o�Q�<�n=F�{��]�̖�=�Ƌk��z�H�I_u�bA��j70����!v���z�����1kk��߼Y��u3��k&�i&�ϼI��sz2�+�)����~��_K�������h{�/�����,<�w�����J���I��9D�
{2��hS��R��ų 5$�?��T�}���6��-/�ڹ��Z7 _��߯h�40k>В�jȎUN�lQ�Qy��p��Qyr�3�%�	�hV��$F��V�~��;B�B�k<�6�ô�u�'��f�.QQ�c����\�������Sp۫a����a홹J�D͇q�]bc瘟}ެ��ᘝx�)׆�1d����}7d��A1B���>]r�OC�LPK�[�]���ljL���8�rya�f�՟�(����5(²q���8�zz�m+Zpf;rJG�k��1S��M��歐�A�� ��{�{�Q�3Z\ǅ�rY���<�*E��!�/��[J�FSId�!#��E��WԔ���g��u��; �@�B�J�[��ޢh��t�F�^*�f_��P�w&T�8�m��g�t_Pj�������v�ƣ�
9����mg���"�Dsє����c������?�,3��z"-���M���5�0�L#n�HhC��PWDei�g�'�)����U�W�!��(s�N��#��/t����l��1x5؞�����:�O
D��
� ��<�;w�P�ZV���Ƀ1������j�MAֵ�u�ϷO��n��.3Q��.�:�r<�S�:��V�6]�Wy���%�E[~��]��M傸<KbNY�oD��f��X���qyﾦ�E���3n��OYU_�J���R�A%�Z����H�����ݶ�w�L�� &��v@�~`,}i{��%��d���9��.T�;}�ǝ8y����pM����v�$ź���ղ>��L��*��>�HEj12�H�@��5�f��+�z*�S9���ݎY��1;��B�{O✮ $t��ݯ�@����M�^O�HI��ch�Dp[�O	�
*i��T8����@8�_d�e(����&ƙM�a�Q�ߝ ���)[svhq@�����(��N�b0Go��H�[�T;FN΁]�����])О�6�a�d�2!~�HܵդPg����'�o��B���/��e���~A6�im��eM ���R}k\ �=!��y�k1�Y�YF�Z����s�pH"ݒ ��֜���5�9j�˝�/��G�lF��ZB}��\�[N�=����^zM3�>I$Y�C���w���sۖ�=X��ut�\���J�E�R�~=.p��ͻ +z�<2�E_	E0ð�lgo��;\2����ȁ\W5��0Xثt�c�_ܰ�ت �F/�$�?5G hk�h�.�%�Ed��@2P������P����)�~���J����3)�k��j�l�b�Yq3CXU(S���h��f��6@��*N	��{��!�6PU;9]:��YѶ���TƝFt.5�����{��o��w$0�37�/��� ����M=�Za�{I�T�@!�z�����5|�D������쐂���n;���+~ߥ���¸��-._M'ӛ�[f�,q>N�\Qo6���Mb�<�,��T�D����KF�N��ߌ��(���`7��*4�I[C��.�ݧr�@��������=2q�-�1�eW6���QM�fD���ڀ�H�p�"S>���F8]�m��6�Y�LD�ʒ�d3�[����6BW����2j�t�?$�c^=��콅]�����*|�܄��G:Y0�x�l;B�]��S���R샟iƦIMqޒ��jf�!@1�2�� 3ۊ�$��p�O⵶�c7�	��BYw����f�$BB�u6N���;Z��@� �Sqf5�L`*HZg@AR�m��'4p�GLe(p��c~����΄ܶ�u�	�f�q�:�����q`�?jB���Ч����mw�\����c᱀u��gֽ��ȱ��n!!v�L1���S���؉����:�F0E������m��E@K*���\F�,�²�`�7�
,��gk%�Pc����Cc��*�P<�Q]��@lɕ�}A�p�βcg�Q�����x/�,��(��I���f @�dj �ۇ�v����vJ������b�;�q��ooA?��=����`�-T�^ͻ��<�Z{-+=:�O�Q ���^�rS�	V������?5�����Ų!���{��Մ_����L2��A�c_b/ۢ���Ϣ�9�hi	\�&�]�ɽ�ʝ��m��%j:��Drq3t�T�t�$�l���n0n��پ���i����bLh�ʚ������IӴ�8����� .تBrޗ����}��r�$ES�
'?�9ə(5>"�V�����}�W5Ơ�I���x���0 ��1/ޱ���?����}��$�p�^Z�x�1��А��Xau����|����Ȉ)3��䃕�8M5�ؘ��W�[/{s7�7�2�o�A:���9ġ��ۛ�)Rn#�F�@.�����-���je�} ܖ��0����"�=�ӌK& p��lk�H�fÊ� �n`�p�k��sU�N-�"��a����u����J�Dy���qN���}e/��-Q�s��E�e������AI>�E��5ot�����'[�#Gt ��ڙ ��/����x@ˆM�0��Ҧ���
�����8}
FY�$�(5���YS$��k��*o �������Wh_sK���
�
1f�ǽ&.�����6%�!n��̞ 
c҇�⦡[/��}�r�t��l=V��.,_ @1�a���1p�'.�Mj����Ế�`�?KWy��!z�`�у���!�Kt�������|�gH�4H��g���s������"C>�\rma��w�5�dί�o$u�V�2o��Cq&7�$B ����	��`"��b���t�Ue��}y���p��0�UW�8�{A��̭�_��&�I�ΐ�,1s�]�i����"���tS4�E4��>,�[qv)W@X@�7�F�B�dؿ�t녆-�Po�/������Vt���t�Wj�����xe�6��y���I( ��w\��F&�u�lن8q�Ջ���[�
+���a�<1����{��9�)p�(}c���[�3Q���Y�-I[�NH[Z^S����`�ɷ����!���^)A���W
����As�
��JA6�����B&���>�i����(N����;ot:e(��dG���P�D~3�9{2P���y��i(�����3���Z^Y�{y�������V�x�9����p������6-��f9 <d��g�E��t�-,��^ź*�L����cJ��-/�n`�7R�!����j P?�(?�ח�d t5�hF�%��B;ER�DE�.��D��!�����̦��Jz^|�m���9���?GR5�vb+`*,���xQ��653�<i|d�&���;$�P�w\a��89��ˠ�8	%n��q�Pb�X܃U~���`��9�M=
����F<ɤ{ �L
�e���K"�>c<�hN"���[�ƽW����g&��K�N�^Y��"�)�4����c���?��/��A�\N]�4m0�n�s��w�����\ 5�GD�
�� ��4g�ݴ$<G�OU�}���P �j>����\X%S	�]���Ԟ���j%�C+�w�X���d��k��>�K�~]u[���)��*�T0&T�^1n��*���Юmo]��.~���9�]�����A��ml��r;�!IM�g���������W�L��qI�u���P(���"�kv�U��T�#��C��n�����5o�>N�@�T��Է?����r������v���L��ʪ��w���f@��u�[�'��S�d'W�Q��f����XߋeO������#�fQ:0:���7 �#�B����������H*�fF,��7����k#
2.���5_�����S˽�����uцh� ��,uF��2�X� � �Ŗ�����fKO��P�̄��)*Sg����5_A:�(����
���W��]���͖���)�j�:ȓ�!ɱ��E��6J��� !E>�fOq
�[���<q�_��~����~���a�o���a"5^E�W�L~���Z��|��M%3�|i��VX���1�;���V�	E����Xh]��.!SP�s�� {k��g�{������l_'��0)xT����������O$̑~�${90�m�]>����kje��v��FNK��9 k;��S5h�VF0���D�K&�V�ށTfV�S��j���Yk����ݾ>CA§����8���'}N��gZii;.z�VٙfW�ޒ�#�w�c8-h�J�e��/����pV�m�L]6����rQ�>!mλ���L+�+��5M�>�z�S�ݽ,�� ��ϒ_Eв��6]�X�L��4$�R8��J�J���{���kG�4��DlP!}8�4�
a��y���*�#a�q z���Ь���)�����ju[C���6˶p�|�a�.�c����6ͪ��!T��Vj������P#~3�\��c�Zm�i��8_�u���$>�uUGP���Ȇs�גlO	���!�2�cL�+DY��ֳE4�P�Q(�Z�e�z�r �o��7���J�O�[߇��:>2Х�B�"�fκ�����xA3.p����Q�<s��*}»�X���!7�O}��k��9IJ�I~L�9S�P�U���[.�#4m���@���x
�q��&���4��}�#XWCa��7�@~_�b�n�HB*-�s�Q>�����жa�]v�]$d������qD2D>� �׬Z�	ٱ �e��R��8fx����9|�d�9�h����Ne�����˧'epN!�t�w���5"�"�|wfi�O��o�łLf�g?i��zFHTuWp��zܠJ���4���F4%լ��\ñ�}9�J��K:�r�(4/�˙X�nVY�:��'�.�deTD��)����d�q7-cl8}`ټ�-q�RN;�!w��Q�Cq���!��(���L�d�Й���:�qiH+�T�X^��q�{2u���AÞ� ��Øŉ�[�r&���M5Zj����؊�y,��K:��˟ ^�PCK`�C\�j5�'߇m�y�ښ����"� �$N�4�Jg�N9�*(��fM�� �m%��{X�����x	������(�@��s80������e����6.�>�/��nnLU�؛ �e�EZ4`��Ho^Z&J|����ފ&,a3ǠF"+�!C�P�	�%��̛�T�J��±qOK�ƻO�u�z`���v�S�$�ӈ6eg���U�{HE�L�(���q�TH�ֱ�=�%�i\�g�#�zsS!��cL�	�ʭ$��\�ia����h����qoQ�R����[��]Lt���~��e��,4�]2���:X�����m��,�ͥ�FAڔ�-���쬽fk�z����R8?��t䥂eT�[*n�{��U�)�Tt[��j��"k[x&Q	�P�ҲʚKg`�h�!���7FF��B���0U�V���`Gȸϰ�����+��/c�;�a����{ ��T�@�@p��y�:�0/�P �ۊ����T�Hn����*@�j�l�_���2�+r�|�å����lT�T@N^�������0�-��#PoJ��RFT0z���A�dq��N����4��k��)ѐ$01/�hN�}	'�H��Z|�-|vp/{��6Tb>�a���זu���
z%�W�N��La��ҌF@��|��F�_�pg�p�m'锻`��S�4.��2S��Q�Tx�Z��G����Z(�ݬ�6-8���%�u��9��R��GJ2vm���&9L~�k[�������I&����L�]�6ƷB�F���etp���l�@Q�߮��
�jo4�UdM=���~^�_C���>���F�{.v�M)��!��,q�qR���/-�D�87��V���h�1����];�6'(Z�)>-w��������QVN��5��jyTx��^5��5t�V�BN$31��"q�C#��L.���o���!A�>��up
��^jg�N�#\v�N���M�[���[�wkc�!�|�[�
M���^2�����oSl�M�K&��Z���2��b�0�8�{u��Pߕvx�(���aґ3e�Y���G]�8
Ax�q�|�?),��8 �߫���7�q���9ӁȚ��'�X��::�f��.-�,�#���X��`�����Dԥ�\5r�y&l�������&/�/��yQ���&<K��WfH\��y_ERO��o0��u��y��r�m�q�O��:�i��/(�n�
��]e��ܵ���<����5XaG�����us͏YF'����@Z��D�0�����/M<|�H�g5�;���~
��D�ESt!�m���*� or�
���h} ң���v��>�l+�&Ӑ�>���yN���Fϲ��� b���3�k��j��vɵN�9���v�B���8*�I=xc�?�V�g̨��)�*P��9�R�_d�2��(���C}`��2N]	�5؆��&����~	���P�U��S[�'�����yz�uWgM6�!J�ɖ�z�:H�8Ņx����brb8:Շ��u�-�L{\�k��f����R rQA7�!+�'��R�����H:܉�ֺ����Jk���`'�#��t4)7hiE��;��/\����������y:S�L�R�g��i�8����_���"+���=ƷaV%�)���ƉI�u�d��2���X� �lHsX�D�zt�	��H�ѳf�66z���H�U�/�������˩}Q����-��t�&��B�$B�������YGcG�2&�Q�xS�L������������;.�U|wY�±�(�6 �qK�H����˒Upx�ͮŇ��;�(���O���\uw�g��b���.O�D�Au@�`��0	' �K������L���K�t�~�^����n����0k߸�LʳKA�� cg2��������Z�J�?�)8q<-�@e��ת!�/�E~E"`�Φz��'�b�Er.A�ι�4,7we*$v@L^O�I`�ŉ���T��.�uԗ�^C�Cn�":"!��j�L����5�QT��A�*�*��U2�tyH�he�57;�b��gB!Ej.wΠ�¦��G(m�g��|���m	#�+�p���xz�f�)��!ö����*z9�D��͂8ɽ�mt�F��$��V ����䇴l]Ȣ�]�1_O��^��T�<`o��<���&Q�d�j&�����;w2��֍O�v,BO?��D�x�7�y!(H4�C��kNV�h@�= ����F�!��8�8Q4B����̒��;��NP�6��sN��jT�X��9�u�9e��ع��J<�;&�������}n����u��k �+�x��j��s�h�����O�I�L�UE���u��Z���v�s�c�������ΨA/"��ӿ�ڰ�6eП�N`Hc�()>xbFQD=��
�7L�\x{�$X����/��K�NZ��>�(_�l D5r�I��M}�9�d�}�X�g+$^�!0�PW�
��Q�l�����cF�/�,.)�tJ|��M�?;~S(�����2�Q�Ȟ�5�b�����'G�[����%?CCD\��B|[BRX�C7�GR�ř�l�ģ^��O�p��*Mˬ�?�7����܅Rݬ�Z��FL}�E� ǠB2"+��;�jڸǲ�~X��u��FE��`�N�̨���S"�;�2rCe?`
�I@�c�N����8AB�1�����K?���-o�����RU_Ώ��i�!�^�B�~]��B$)L�a�5����)�!�e�Nd{�-�]�Oå"J�<{����2��9�� N�h�H�<�~Ջ[bp+`�k]��L�Ж2[]��	T�h�#�K21	>X��|?� li� u���z�UM����U����3޷yma�1�\.�"���Ye~����z>r��Z��X��k�9������W�$��U��N�-K�#�р���cAU�Qyڪ��:��#��APt1���rų�;� A�_-i�Ȯ(�C������v�09{�*��#�D��r+��-e��#!�7ۼ|��Q`p�ƫO�`tN�6�*���C��T7"�[��(h�
�ꞎ?����9�7pG��No'�#�?S	sMtJ�Δ�*�y�
�t��Ô��p���޸�����Dص�;sn���֔|�T6���@X�/�+��z�Y�� �^ڍ���9q^
�(���tϵ9�KT�B�e͸N[=	��l6�� �Ju:bn���@�:<��[Ħ?�x���:$�����ɬ x��u�)oG?l�_��@�t�ě}f�lz�UM"�zL�.�aW䵓8�������B��H�c9�������5`L`�ԣo���Z/����M����r��)O�������Ի��%�,�~9���t�*Y�j�~BQ��2xO����C5}w��i\�Lo�t_���M������|�f��1	i�ϫ��ߢ(���25�����s����^�T����Aln�b�)�>��R�_r�?��\�7BgJ�kԣw4zPE:W�.�^�W��15n��妀DF������o3Gi�P^&���	�a�PMb`��$k�i��+3�ɻ��t�d�g��:[[ıg����G��� [6��	c���{^44W�N�M7�i2��p#������p������:�����*ip���Ɂ�0�Q�T23�S����ܛ�N�|9dP�Q�q���:jܕ��[&Ɏ2W��q�2�xd�j�b��rL��i�;;Ż�]�~��21(X<����r�$�[g�Ӂ�(�eQB��˷Dk0�M�E����\��lp��PD;��2�ߥ}���~Oꪹ8՚(c��ϟ��A���aT���S�q,ӓR�+�X��<�g�I��/��)ah�}�,_�����i2 ��*߷i&v� �����3�ީ�:�X��-�2Cqj+>B����ʘ<F�1Ȅ��RCt����xQw0�SZ�xZ���s<e�r���(�d���g,��U��tT.V�~J^InQcÇ�ǯ���:�=T;cָ��x^����p�g���q���4��W���4תl����}Jy���}�5z��i��FIz�fO֤��ń�
�a͊#��U�0a��|ќ�s����,0R�SE����`���[%�d;�-z0ƶ����
��Tp�T�M3���� ��E��
�<��)'�g������ԁ=�=
��|å�Uo7�-�(^ɣ���؀�'h�ܮ+^G��:�j7��@��?_���H�q^�Fm�޸>q���֜z�y�6*��|�D{A �9��.c ��](���5���h�޹��DD1�1KN%����K����p���H�_��_e�ؗ�z.���;
�iUV�n\0���>�.�s?Cf���\�KxT����x�$ux�TJ;�`�I��S#��{f�H��D��ɹ`}�\��u�{�I��I2��k3(���=;*��*���3�f�2��V�8׫א�Bz��Y���l6��JRe7�l�Nn��ro�A<�>�s��
�uh��mv���O�^�v�p���D030�x�H�?����P�2[�.�?�+Q�=Y
$�;�
�?�'��
־g\q�K;O.6�-�\>��S`͹.P̥��]�/��Jo��JP��;RW'��O�@��Ly��N�qj#�i�<�y�٢Г�̺w-�z0�y��pP^����%pG,�y��g�%M��bR)�A�F������Gs:gxmE�U�`:I��K�)N!;���7��P���\�˕Cʾ?m*�wV�=E/A�&=��YI�H�U�3&O��{V�"�Mw��q�էx�2�In�AZ���^���T��7j�o,n
�Q�s�R
�i<���v}z"KzM�g����$=9|9�e6���H���8{*����5�	��͌bv�j3k�
K��8�̤�9
=�t���C+Y^̬�[�+�����UpDI$����В�Q��[ȴy?ƹ�m��<8'�����75�O�%�BJ�M1E$���?��m$��+o\!|K���:��`@Z��u!���%|����c[�
���|���X.P�J$�r���Ay���zi�rKY�J�G��)KY�()�1(U"a��:�E	c��M�O��u����2�3Z�O�F֪5_��3D'����M��4�X�����3�̰�;���c�Sl�©-,Jwy}c�k*2S��T���$��$�w�$�@(5���"��9"��eZt���z $��5��tA�қH'�./R���SF3�3`k��f���8��|el{B���������n�2�s����ӛm,yՃ�k���)Ϋ^�.�}t�*_�U)�8!���ژ;�@�	\N��հ*%��G�}E����\d��Z��˥d����柀�!��7�e��)�:��m�vWi=���"���
��u�0�\�����it�&/x�S!�RZ����|`�O�D&�E�|-6pK#�.t�'����E3r�jO�Eǣ�K$�*�QK���Ȣ��< ..פ(*.z�g��&��M�B��F��;�~�r*q��	k֊$��w�bSJ�F��c����4#����o�'����T�݄�<:x���3w8���N#r�
}�������u�;�:���w��Q.)d���zɺRc�B](�T?h~�nI� o�m�S���2�%V�x�P&eY�w��g$W� ������s~r����{��с�e5�^�*s�J���!��Eh#�	t�gb�p���l��`IO�Ȉ/7��s��L�O�B^��Ml���|��_�S>��Q��r���d���~i��
�2��ӍF������ |������ ����/���8�:�JƌP`�z�\5�ѭ�Yo�cD�lހ?jCf<r���
��z�N��6Rhǲ݀z�/��O;�B��7�zE��5��G{E�y��s��[��l�sC3m����#e]�#���%+�8�� �y����ː���W��W�(b��)�ۨ��U�a{�S������v2�i޵r� �?^W�����!�.�<��7�Q@8�˼����ܙ'�쇰�!��3/k01����-�������UFմM�L�+�g`?Y:�=EQ���v�2U��(r>�C��c���}�i�N5Mn*T�=�##|
ݐԀI�`b'<�F�s뀨4;֟�达���>9N4܉�>u�~�2�)o��l��q�j�6-**[��8�e��噽O���H��#�z^���z�>�9��i#\���7~'���f�f��6|��@ MĤ`�99����Y�^9�L܅�/.=Qb��h�n�n�#@O���G4=�p_A�iV
m�3|,Y^��A۸�S�0�K^�����䒚����+�'qW�.������%�ިe��}nބ��=�<�Z���n��S`����B�G�Rd}⩣��I��/'a
'߹hT�.�`�X:B@"tW*���/��_��ͦ8.���ґ7H��8���]�4I��]Y�}�F:�i����r}1;�.�{޽�ȞѴ�|� c����;r��/�׳ag���A��/��dʘG$�o*a�`��gɵ����@�篠�j'x`ς�0O�k���j�ܱ�V���cץ��ޚ�������t����ԾAc&J�@����i˳��)@况㖊�E�n�����T��N�nК��+`���P#���������M��n�ߢa���
#JR�q�yU
u���b�%Q|>��=S����
[K��-ׯ��ͭ�i��B��\�B��7�=JT'K�7����ԩ��e@R�w�0ܯl�1�`���ONt�&vq�#��*6
�3V�u���<U���aչQ�s�8��,9�Q>��(�B��4<:ب�}�l p��==l�J7s���;	���ҝj܆�M6�� 4J�*����J�����X�\YV2ǵ�/�(Ƭ����\��� ��Xt�G}��78�ʿ��0t�a,D�d��W9�;�p$��\]y�����>��.��g�j�B˨+��*�5	d�t����G��zM�V�J�h7��v\�$o/�s�R{�M}�6�&�@(ȃշz���i�Qo��?��<�;��vzԑe���Z��R��*Б%�,4�*�h����רZ%L�*w�bG�@�2�K���T�T�.kկ{��v�r�'۬M$^D�f�PER�p�s��5�+��6�����ۿ�9< �sG��n�@�/���y.j	zc��a�f �K��$@9��#�T��˃g�+ ��`l �ĺ̪���\��2Yˇ���#�O�^��6Z'�?�(��fXR�#�0Y7K<�4�`�:V�P�AR�a�<D  ]�[e��f�;��s�ny��1+�m|9=WO�N�}Hk�2�[���D�f@ \�i�5� ��ͮD�!���o��y���{	�݇�^��&��<ɺ�v��VA��̡3g�%�d�Z�3�e:r����l�[{���X]���U:?�D��p#�f�?���.�K}��Fu�pI��7k�ٔJ6��~�\z5���8�ヾ�^Śm�V�aW*HXE�{�=3QWك�f���rzcw��9\����Վ���*��#�D���⌑�MW����Du��j��W��IHmF�|���U.��I������W��y��[�M��H>#&D3�VnY�or�������)�.��M]����A욃e\C��E����W�:Yꃹ�e�[,}����T,
���ap�Ӿ*�v�R]Bx~�3N�}`�q��a�4坎�W77���j��:��'`߰��{l]�����6�K��B�<�*wtu�jS�O�g�ɩ��v��m��}�'��y'h;͟����.��*T�ZJ,������f���ޒ,p��"���VМq�ڹg���)��,v!�Ż I�ʼU/��/��u���lB�oȖ�,Iv����t��n�����}��0	�m�A	��ߊ��Rg6�!'�� \�lU�NZ�	�skK��^�V���I�jI�ѼI�ʛ��I��I�#P����X�P�\�_
顭޽����Kgzk7_!�0�{�ڤ�c���������p@qO�ԫ�1�E�z�L>œa����v?Ja(7�m2�$[� }�1Ǽԡ�Oq{�Os)�ٹ��9��ǡ։������?�T��[�^d1t���$�3�,�(N��V�=�@F���[��4�a�lT*�0��t?Ｄ�W��NuXi8�U�0���<����&jN��Bz6-�-߲�A�7.��5�Sa��h_㛒 �fdp�2i��F8���{'����3�׺;zIP��?q�ي���8�}&�#��qWI�w�������Ա����/��^qڄ����tν���T2��[�m�j��T+FĹ9�t���PҊ�����J3#K�F�0t�A�XF$MBy�5J\&��jLU�t�n"�儦�1�����p��k2�_� �؈�k^@���t@�6ٵW��R�H`S���`D���}t��׳:��b��t��@��Xʭ���ݢi$7�:�ˑ�ܥ��.˘o�ˮ� �l�4��bе/m]���2�rNL�X�܄Z*>�1�Vf�;�Q(t`��k��w���)����,7��sm�А1$e�`g� ~���`�.Hp��p�����(��ɋR�)	2u�"HҬ�:�Ɩp<���a�&�ۮt��s�G�Y�Y��H����-� ��c��Q�l�����:�$�ߙ���[��
��WԒ]N��0ңp�%�꘤�'�$jj��,��v�U,�͸�$�����t*��N*��hE�m���R~yzi(��ہ��U��n,� ���p�rV��pk�iHY��_�O9-{��NbJ��vS�]�r~+��Y�P�/b����U`Ȩl�9i48�lwW�{^�#�5RJؤ�	��B���&��!����Y���[�}?3������J����b����Z���9q��ͤ��*�r&�<�|9��]z�G��J)��`�!����5���&苶����h��4�j	�8}<���pM�/���e
]E��K��y2���Ic�{�L� 5G����XU���S�Rv"�Ik�3�����j(y�������O~a{}����e9�r�)s�!K��1����h=_�ʛ�<�����少���st�2�ʿ�}^��|�}	�%ax)�3�ge��)O��rC�IX��"Gw�]���Ǯ9�e���m��di8�rb���{M������.�3Ǔ�i.�A����z�e�o�F�%�dN�Ɋ���s��w�O��di: j�gz��P�_P^I\%�m|_�u��L@�0�Y}4���{>e�Q����{-j��$��30��a�I�Z�0�KtOP�~¾»T�3�Ð�36�k]Dn,���Sы��+>�q�V�?Vfrp�����W��i�@�oɣ�(�%~���c�[v��+4�����-KI������ɰz"0cN���Ø���1&�}����r�g?��e�dL�;g�K����<d�]tA4~�������NFQ��A9��m�7�x- ��R�Y4�qZ�-]��ڙ)k4��Xg����r���>�\��7?[�[Y82U0��ދ�,�3e��xEN�� ���*�٭vFp��V�Nb�X����g=���Y��#(���[�]��	���߷r@�w� TL�m�y?E�B���K!������x�Q�1X����G�Q�4P��\�6�)K��E�������їA��U�6&��fxW��?2�b.*x:اu��q�~W���k��V��sB����)1��ۃ�!�!Zn{�8��	���|��! PҸފ�m8]ڳ�3M�%z����� ���S����� /v�U���u���\OX$��,=�L)ѳ����wT�i�K�}S�Ҟ~y��ģ�^<d'r$����7����#��׎�G�}Ӈ���债>�h����<�a�^bH"�>:�M��D�8�C�i��O!0��jc�ш2�Q�y��ܰg���9�W?j�~u��W��v�oɩ�ύ��؀[��ҕ3�4�٭E��X���,f}Ăf(�a�LDˉf��ސIّ09��s�Eq��nб�W�lǅ����G (f�����=��q�,y�"��.HO�c+��Q9G�L�4L������'�9��K�d$����\@�;���1l��`|��xIɪzVxğ)�p�g�Q���nvw��U�z���Kn+5��\y�]d�z)B#�wfh�1w(�����S���亊��5�D �[��.]fzQ~�����=����0�g^�hJ��/��^%�L\����@���\���W��ޓW���u�[�d�v$�yY���<���f�h�v^���{�]�Ҁ+�@��t���ÏU<��y�e�?K2QqD<�xK"E���84���|h� 0a��
&8��N~�������8��P�Ŋ�U�(Dg����X��c�΋Γ�,"Yl�j���h���K`]�7�f�Vl�������Λ->(5v�{�B��S_GĠq��0�[�x4gdO���yN��(�{�P=ț��Pb��$Aه�~���m	zqn�=;%F��fd�J�[�u��O
b>�j�6��S�
d.Bi��=�V�Lǹ��7�KI��m�>��
[¯��%L���t�$t���2�I;�.�b%�I�Ҁ���[Jϖi���a��kJg�O�A/��N�o�M˟���v6�Q����H�=D�)�������6�q�����Vao]��~����R{Z+�ƭ�5z�LI�sKЗ����݂0j��ud۴�Pح��]�����b� �W�R���m��w��De����(� ��:�ks$~" GԒ/��aLĒ���]3�4.Vm�b1�������Y����D�,�x���`Oő�ϖw�b�zQ	�yh$����~Ғ�u���$��[qb���>��{:��+{�	ܝ���b���W-f�V�hzӔ�Y��b��?M�[/# ��3q��8po;��=���j������`��Z��� �#:����q홾�Ƒeb���v��ۢ�|���Z��6���2�`^�B1V0Zi#�N�T'�luHY�4�nE�{�I)..��Kl�j %���Y�S��57Cxo��L�d�h�E�W��T���Iw�>���%� �%E��8�G���,��`ﵬ�t���U~:�f���}X�������C~(�J銕�@Ԕ���w��/I�Ny���=�v�>���I�l�K�Hオ����/.������&��8��"0~(�<��p5�<���8|�F�"��;��"�����h?�0�rգ��_�9Q��%,�x ^��>Tq����ں���Aj�rGl� 
F�
օPZwT�,C�ť�=��2�����ىo��e�r��`���-�X{���{G��]�?����5C5%Us7�j;�.?e������� UP:��7�r% pvˍ�w�q��"j��Nˠ�P%���/l�4�Rk�}&��Rs�T��i�u�"ciK�(n��3"Z�ufC���Nl�f=LK@i]tm����Wvϛ��� ��YZ��l��/GdFk߸G�q
|F�E�����
��NJ��v%D�D�4�)f��s|=�@�3�=�rk쒸�@�}���e�;rTʁ�!�E�<P��ޕ��M�Gau��y�r�h1�r(�s"JvYc���_�[x ���yp�$d�A$�J�w V:@��8���{B�,�=�p��Ln�hSkUa�����P��`�~坼;�,T[�Jw		^:�*�����v��Ǭ��z�E�,PCH�g�Ȁ�y����Y�2=
E�&`Y��k �-C�#?�ޓʠbw�d���#*���7C��Rٝk�[�Gm�Jƣ�� p�C�n�Χt��0ty��M�m��\���/2�˩Y�l�9���ٲ�AK�\9G�(P�t�v�� �EeF5EGK2���q@~ed$�{����J���bAs~:�a�OT7Z��8���K�Efvo��g�n@p�Wy��y�{e6�u͵j��yn�{��ƛ��~Bj��%�K
�,�Hw��0� Fڍ��A�������=��n�����^���WU=R)����.��D�g���[�}J�F�ʻ��s_'3Q��p�*�d�����5I�.A�,=�@����B<�Yѣ� �Ή��H�[G	d���|�œ��x�x�'��ˉ�5��M��@�nDY�S�b5\�'�/�r�Af��!��2�q�=-N\A�����<�U�����G�rn��i���DBo�U�祈_0��U�M�7� k��vݣ�3�Q��VQ��!�Զ������.�R.���:����tAn:_�}��p�s�yY�K����.�R�kj01W�J�r�sqؤ��S���2��	�"�OYC7u�t��#�-��'�����3�R?��hz���-��U�+�^M�dXCy��u|=��� ��䮅/���a���
7���0o��x)�
i^�(F�K�zeY^;������������<�?���g��#ס;K`̗^z�D��B���&�
z,�\$3�x�e���U {`�/H�.MP3�]�q�K����Z��|�Lx����d�| MO~���BO�6-Z����GxK�3�4�]Z��ZF'9	^�69<�+�%�Er? P��Y�$t�ZE%��W�z����g�]���R�m�Eg3R$d /�j�Y,~���( 1�S���(6�:huC��~�	���'�H�Y[0�y��r����L�>�D� �3�<����p%���s֋:?Y�+
��n.Ԁ9�v6ބ(׏�zB3�p���vj
X���#�d:�`&�e�O�ġC��
m������g0������l�rvQP�{9��1�I-.d�0*Y����M5��V�3	�\��0#�\7�b& ��	�2ۣ�A1yR&l;,��$��%�����A��V�Jvȍ-��jZ^�?�lmov���25=[�wū��{犗5�kt�(f8��袻������9ds6>4��5 [���߬M=5�L0�[��2�Qe@�D��E΂aKȣ���:���ɖT.��ݒ�Ƃz����gw���3榵<p6�������I�<�8լ���;U����9%==%&����kgS�!}���`v�o"$C�Q�9�/u�c4���L_㤘�qR��?}1����D�u�b�Y�I�ۮ-Ne�国�։-m��e?StR˾��)=<�-�:������;�Z]I�l"s�tʆ$�녖���p=e���=����k-����(���=��u&������̷��Z���)�$��K�A֯�1����%����6����J��g���(�]���r'J�����"�4P��#Q�ڑ��\����2��=���a:�xT;,�!i�l�3�"��_�.5�0Hzw?%uĐ��u�1��Ǜ���s1����?#��O�L٭��G3�������8�g���|;Q��n���L�ugS��v*�.9�v�Zs����dý�����魫Cީ6+�FmI0��\�����Ucv:#��(�h1���m�g�	k	'�vM��_�� �Р����Fp�-8����B�;v5� ��wb<��lß�Ӳl�q�EA���{ToKlep�)�����E������~��W�s��� �o����#�῎K�{]jn��1�"	���QC��,� i�����:���y6�id�٪�m�+N���t��N��Y��s����n�G�<�ċ���-�{����p�ڑa+k�*v8�]t>�m�@v�͊��U1�+�D'�F�"��/�u�6h����%�e%!^��^� o��|����R�p���.fù����1�5���(>l߶d]��VQ����M�[����\�ߌ���o�E�uI�g�=+L:<|A8�a��w2�v�����!>���{j����?)��>��ώ|f�N�X����g��B�N�1N�c��G���F�]�f%�̚aM����b��W�Ӭ��ѹ�]���&d����d����ɵz������ȮIX�mYt������bE*�9~ޤ��.�L�&������_�X�P} ��*)�� ���!��o��86b��H$��C������V�be��A:���S�+�fS��A��b�S�'P����5��y�8��V�Dk��� �*��S�@Y�L?,�;����rYCMd&���-�mzw�s��n?���C�ڎ|���FW�(C(�,��4.���TH�^gI��%����|@)� 3� �yU@U%d�[*�Z�s�^��/85+v����������C�J�2|�R�6<e ��Ia��e�G�0�A�ϯ�h�2�����~�%6�}IC?],�}��o�<�%�����6w,������� ���0Q�A%g��V�w;Ђ���h|����%s�QY���Z[��=z��Qj�������Q;#�3��N�Ӆ����N�ύn�q`�3kN���8�n�BX5�B5k;�'���bw'�
��+��7A�K��1�&dU����@9�w��cl���;	$bO�#n�Χ��g)�'��z��۬�	/Z�yn�8��#�5Gx���4	�$N����s�x���xf�tx���(�ò(�*�-�y@i�w$�v5 mo�(#� G:��|-Cl��';�ԣdPm:��LXn�T)�0�SY����~n�Lv=���~hւ=�zg ��(�j���>cY�z*�B�,���]�)��%!��^�?�G����$�ߝ;F��f�7ͧAB6��P>4ä ���`ȋ��>*���OZ�Y.�[k#����66\2��^�b	�.ֱ�-�p�EV�Ƥ�p���ՉT�x����'l�E�<i��2�$G4x�;f $�蛾Z�b,� m9eJU��6`��i�ת�%-��Dyg�x.f�Ry����D�&n���py�����������˗�w�������d����i�tM8#� jO�㛝}W{G�����H�9�!s6�����p�
anB�>��n��7�t ��>_������,�߃$��3>�b��ھ�ӈ�P.�֟ꦏ���ࠫ��.`���I����O�m�K�5��11G�K�v���7^CV~{dA��b���{ Y���Ege���BS!qo=�`�\��P|�5]�iE)M�L��x��S5ā�zTO�4���{H{������t����8�~�Y͹QvE��,�*��X�ȍL�C_�,c�Zʲ�gLoa�x�2zM��'�Uy�5��m����]}�p�!�28Zd��Eh�,T��N�>�찥��\" ��p�(��G�A��	���͝�g�R��\g�ڔ�����g"lf�j&M�{)�u���<'ah�D�9�OP�=RٷNA��s|,bh�bc]�A|#��F�%��_���{k�;��"�'5��a�����\iL�/�-��C��,DQC����c.���^Y����1���I��`�]��h٨r6Yz��Ъ]�=�MŻ#�ZIG���h������{��D�]���e�����t#�5)��~��vU���DI23�-�״(��>�PS:�i-1���نQ�Q��)d6^ms�IX�&�a��xOIlu/M�0dD�R�k,&M�,
c��z�aר���ѩ'7 S��ИU/�:�<��揞u�G�BRiqN�hQ�dw�P���v�oe��vY��:"!�9�.k�J��V�ہ�8�h����9)Q�Zz��4*�c[�M��U�;�ĕܡqq���ݠ�b}���TP��eU�����i;۷���&c�8���#��U&�#a�ٷ�!�>st��� �aҵ�u�;��[��Lލ����]��фR���X�e�H��=�~V9�&�+Ӭ�m]�C��9�n�[��/��;dQn���X$���
�'*�8�T�-���t��u�����+(��_%�r�qRK����~�9��Kė=`�����~yP��&[���5��c�;�?r:L#f)�w�.Wa���J�68�d# &\����'z�ڡ;l�ܿQ�=�y��o�i��WTPC�u'dۄJ����r^`��Ҿ]rs�����I�}h�e6h���6���7q��SL�Pܓ7jlE���\�����%ܾK^�S�IwZ���m�ٰ�a�o핮-g��]���1���{�i��=��Y��`�ks�[B��yr���v U�����:2��N�)8+�`�uE\yk��6�O6Eƨb�Jf	�P7��r/�}�-�}T'�G��~&f�Y�I���
�z;��<���`\pCi�`K�M�wt����
��;'���,�~�)�_�L��i�)��P+����0󕚯��pJI=#c#�d��Q6�F~b]��� ���I��[/�Sh�Yv�(k흙%V��l�[K��Ǿ6�a� ��ٻj�^Ś_~fk6���^+gmU�{?k�tVŸ�����*=,����-����8��kȲ�غ��0Y*�u)�!@���Nd���� N��h�K�n�׸�c�����<�Ԩ�D���G�kY0U"0>�h��פ���[Lଽ�<�4O�'��x�B �9v�9�G�S�M��t �h�C7,�A�\�A 3`Q�ґ#E�}�Kj���D�����i�3��t�����Y�8�)�qƔ���>��k�	�4��1ݘ8g,ķ�7�e�Y�8@�+�f����.P�7��x��hچ07r�ꍤ8�y±�bB���R\��\_pzo�d�'I�c�V�d�%�h�1a�7�,�e��_�Ũ)��3|��+1��ə��Wm���3r�S��e%��G�;:_S�
�¹r��f�"d�\z�1�����<�{�x"���5�쭚V{���N*��)w��Xd���+��gv����(	u<����fVt�T� q��Z���:�� ��mŅ�3:���p�d���������	/_�%�ޡ��	��`�w cD6��wX:�Q�4��~~cbu�~� N���^���� ���h��α#���٢uU�V�v=v�|�-���������N����{{D���A<���ୃ
u�4, x�!�}Q����2�4 �g�Zo�eڌ%�BJ�1���{nc�Q/E�1����]~
hjDGU����%Ĵ��%�("(��w�>R,O�n�����:�9��[;�!޽T�Y/� �X*U.�^o�Zc�`;kً��[��������^�>2ߋ��î����-ah�x��ru$˲�C�c;�9�.$r#�j�o�y;ny>J�}�0���Q
3�J`rl��4�F�.���w�O�X�����@��U6ue�;78��j�4��d1����hV�m�+�!���JR$��1�>V�����W��n扌'���u�T���cɈE*e�3�(���u��I�&t�^��=�-�@��&g�d+������SU���K��bv����e�ф��)v��aI���,���3� O�V��>�9w���e��׺�z$��> ����Yr����4�<Y�o�[�iӻ�_��o��t�k��?�+������wQR �Q���λ�Mu��d�Iu(�5��wR�?���q��R��d��^����3A���4�y���� �$%d�x�t7+e�dR��"�	���G|OV��Ĉb&G�0�����z}!8I<a�@\��BW% Lb3p�K�N������:@a`�#�=�֢n��A�b�AvIύ'����ۃ����MNF��̊4+!Y�l��@}�����pq&�q��/~B_V�N;ꖥ�*�+e/�G�<'S�4��A����V=��p�G>���2���"�$��t�|�I�[�C<x�y���;P<��S<g��*��U�i}F�4"���J`�
b@]�T��JnG��Q�O�Υ�� ���,���@��=�79���s��$*x牎�^�����`�d��w�<�ΐ0�ӢQ��W��'O�`A��Dqp]mZ_���l}�Q�q�21,���t�i6��S�O܂e��i�tR<港���B&�5�X��٬��#wz����g?�g��� <\��R���}o�3��u�n=Ȓ�O� |=���v�J��b<cYxe����&a^�_�mZlS�̲�D�}dL?�5�k@0��Fg��!8�ȼ{+o'A$��Q	�o���J��	��A^܉`J�2r�����r17���Ǿd.5�dyid����_Aj���0'S�0UŰͰ�3E\4k�fO�ߍx-�d?�������� 4�U�]�*fh�q)u���1�5#��W(=A����d����?��qV�E¼VUNH#|��U)�4����@X�ox��E�Ln�)�W=r���]>�PlQ���w����6�'�8D�����i�:�[	������SH��8!Xčhb�D�Њ��z<����_p�t�i�?�k2�w�W�Df�}KV�{[ݍ��G���7:�5�Ϧj�{g�����zp$Y�<�
qAF�c��1�R�9=�6|���*�x�3P����9Z����(u��51�ؼ���H��H�*E�>�~�߼SA�7�O��[�ȟP�"�l�=�%��xc����5E�D�MgsH��Iԅ�fB	oX, �l�6ҭ�W�ū-M:g�<�۞
g�O2�1��4D�˥��MZ��`��1t�P���Ԅ5\��6�jv�m�X��v�����xj����p�I�����Pf�� ���iC~k���H��Gá�l|��<�::X+Hj�B�yQ()�c��`@�0	I��|)֢L���,{XQ�f�2�N�O�v�[A�z��#o�lq8��̊��>�T�@�Ep9���t����V�-KS�3`��;���9���w�	�V�aw��`��I��@����|v�2 �~5�����@jt�r?��Q�PU�@����D煳)�g�ǭ'.SS� �B�����>�ja ����32��J�̅���Fl "�	2��,�´+G��#��{*ҖܼT��{z����O�q��,�B��	�v����*������{�^��ݟ�cO��<@5�zGr����:�:����(�����1��im������"LtÆh�Ҁ\.'1hwJj�O&�U��<c�_�ʙ�`AD��z`#0l�a��B��0�ջ��n�8��C|\�_i�N�k2�9�}�OU�NY&L�NMR�^%��X�KU���U��x���k$�������Ot����J�1
�g�x�y*պM5rT j�iN11
q4G'�Y��2��>��;^b���ȿpk�#3"s�m����*��	-�l1[�����g��M$L��Q�7�g2XB{ݰ��8������V�q�,�~O!�� ����d�������>K3� Tƣ�2��5�4r�C����nA�}��O��΍�%���h����b���'��D�)���=�+C�����̅�n&ƫEȞ=QNO/N4`� �%�gJ���m���+�4v��#��h���V�����ĮOq#�ȝcq��"�taZ��&�;vh�]Y�hS+��
M;�뮵���H{�Ce�9��zi�X���	h��,��q�O�ETR�;��n��Ë��d���o��[�ŀ(G$9�.���i�;���:�-* P�βʍ�F}wQ�Bm

��7E��#?�f�Yc�uȠ��|����Ղ�"ў�!h������>{Ϫ�Â�ĘCQ��wH��7�^T�Y����
�FT��*�'|�_��R>�&ߒLƭY�{����9���l�E�]��f�H�=�r,�Q��6��X�H�#C��ub�Un��B�C�������;~N$b��Wg���I����G�) wGG]�JZu�|C�	�܆=�����]��2�:�љ��P_�~4-���J��=4�+2U�g�s�B���o���~�~b�ĩj:nϗh~�-5V�t��k����t�n8ٕ��Y~P�1�V�3�}�C��~�PU�`��7^�O�z��{�3�	Z���n!u,O��K�U�����&�*���v��/!_��ã��j�W��ZqG����Z�K����������K�\i� p�2�^q٪�#g(�]�:���#��)�DS7���a��K���>���]W{P�v`��a >�{�5���iZ!�KXb=�������-]t/'(תf�3r<���R`|en~�E���؂�l�uE�4靻���zAG��6zҟeh�`m��lE��}���͖�똘������7��a�Q��V���|�h�5֣�_��8ڡу��"����������K� ��V�iu�SG��#�?��7�=kƓ���\�PqW��3�b7�dV��n۫8n��:�d��a��χX���J�9�lŶ�'&�oÏ�CR[�����1��ן�-��A��h�!��;c��h}��J��qF~u�'ˁ2{�^��������XB���n��N|�76\�D�`RT7��"�1�*�3zEy�Xùa��f�b���a~�����閯>� ?y�C�a�H�S���k[���i1?g�;��s�+���$��A��W*�(� �;�V�N�+ښ�/i�;r�^q�:}�A������iW�|C���>ë���o�(�W.�T�#�����D�� k,N�����<4��_�e[ZV���85uu"HYrU�}K�!�b �1j�е3�e�N"�ږ$�l(��.st:8�cqR�2Q��Ր�������<����E?	yZ�i�A$�f�;!ȋJ6J�R�#�mb?�t �ʢ0����l�cv����8��ݞ��.�M���	����;�J�2�.Niol�z�&���k�+T��i&�3\�/1��������װg���������6E�+KL�gIBvW�EʦW���nn�)Y��%�Ÿ@�|�=Q�bҭ�*�.�����v�QR{{%�|�1^�hVmFNE���4�O�ٱ>���t�"Y��E���Q��R��AlXs�1-P�N�h),�)������o6�|��D�]	�5cG�֪�s��<��Y���_iҶHr�ҕ{��7�"��=CA�gPX����d� K�	Y�A>�3��ռ@:�W�D�����^YFI�:�?&���G��9�}_�� Bzړ�[_�x�ISR�Ε�Ͼ�	s���_��l��-[������)!���Nx?���DY|�} |������c
V�l��P�ñ�@'�ۆM����l��t��5�Gqb�D�DI�'�(��6��O�P2q�s�r'�TlD�$ ��j@p(&;����q�RCK�td�+�_5 s����l��������� �9@�g6�O�N,���S��S0��iM��>�Udۻ�~"�=�ws-4A���M���կR��y�Ns�[)qt�sa�~�����d���I5
 qH�؈�<�"�dD.9|�A��@�8P�u�}��ly���,����5Θ���?��q�6�S��U�;�S`/#�������+;��(h#���N����s����!Cr�Gz疚Wڒ��Oxg"�0���ܧ�8�@W�\d2���*CVƸ>�$TwV)���x�� ���<WO�4jE��P^@<��)�0 �W)O�]�6��	�%� ���I��(�вƦ}���œu*-�f�7rC���	:ޖ�)�g��P�ArS8�Tz��j��U ��Bvh�U���֋���:ו�fc�fH��u8o	���~�u�)��j"0*�%{a�|�9�#X��+�'��HC;J5	�[��4��{R��/!�����a�_E\�w�����|R�p�Q
��l�K��17`�lu�Õ���E��w�qlnuQ��� ��%�V���M7/��A\�O�S��.���8��E!�J��U��-��&#���A�� ��Z��1�Y�J	�*��p^R=Q#Ȥ�_��Ȫpħ�9�=\O��lT��Òb��#�M���EĹb�W�w2��l�r�ӌ8���L�1�L`�6�N~�h|�ґ(o` �eS�)j�z_2�6.�[B*^�A�ߡ2�\Pt	����<=�4ܐGۘ M.�q�P�U��T�{�2_�ɂE^%��,p��H!q2�"�>ZA:y��_*�P��)g����k�/�H柣x=����xӚ-��w q$"���F����jBwє��� <<������pl�L����̓T:���b��8	��u��u�L����vX���N����Y��o��A��%P룿�"��r��-'��cb_8���v!,/�%W5�L?vAQN���=�{-;�����H����S 6:��!������~��b�
6yߢG�s�Aw�;���"MN/��suFH*�(�oؔ}�|���pK0���VFv�MM��� 8p�]Sz	W�y�{�+Y�c��88���3���6,b?g�Y�Wj1�K-�'�G������y +G#�ژ�
�"q�$�3�oYA��Y;�����(�n���QIN�	-�Oq׿��&0�s-M�����n�'�
����n�����8�2�Te�}!D���͊zi&��<�N�e��e8�!�K{VYOx�lxot�,��a;{�����
�8����\B��)����;��q��C)�u���
��"O��B�����c���^s���ٻeϛS�"�5��?m삋Yv�����i��`%GT��_kh��v����X��,$�i� ٸS�mTMm����g�E�(L�|d�Oip��*:�?�Ĳ@��r:�h@�ǒK�������
�7b��~�(��7M|�'��&ѫ���:%� �Ux����[G>S�^_����׈E]ee2>|}P���C�	'�@Ey��:f?�ꠧ�	Ԋ��j�D�ZG�9�'�O?��`M�}7<NSs:V��qgt�S�$�QW?S�r*��x;�p�
h|Fg��_6.)3��`����E;�V�K��F�P~���)�n�a��_Ϥ)����>lE�n&n�m�ŭ�O.E�nU3N����L��I�?���s9Arү%��C�\4q��t%V�p�Fޱa�/u����(jA���g�b�bII�]v�Q"íU��0l��r%`bR����-�|���d��*�G��,���kA�vS3���&�8�&�)���o�č�x�y��[d�����]9U���C!S�%�PlcˬA�*-�O<�&���C�A���)Ƚ����=a�.t����#�-zެ�jI�&J������O&3(��ϲE��^|���]g�(%g�d.��6��N:[�0��P��m�%�G�s8�٠W{�pd��W��˶.ٙ�h�[��[#�����8��
����|\�'
��TZ�(���3!Z��L�>D���%\^�U?mԾBb��d�Y��0����t�8�*�]Jl&P9���P	�Fmi�qߓ���}?o�ͻd�:��N53�ʠw[Rn7o�����lc��~ylXA,��G7���j�Ń��	�o���+�L�82������N�{p��_G�WE"
�h1ϜA���e�QL$}�p�m��Ԉr@)d�/��`��+��֓4)���*`	'd?��c�H<��Y�+ <�L��}�~��.ݘ�!�ٯ#�A�p��'�D�h��;��㰌�.���	{��y��,�N>˱�e���������f���t�t��c�{����_�V���0���[_�eU���=e�0եc$�� ��ܘ��T 1�1�|6�"a���w[��x�>-�2ʶ��D�<I~�BD�z1Ƌ��sR��-+Qe�kׄN*Uw.a����r���3��T/�c;v�C-jz��.�f�1�����Z�i!f�W�{,-.��T����^)pꒈK���W:�����2��sy�246�?$���lL��T��b�g�(ۀA���o����~�f8��c2nVroy*�����p�����ՄOp��{��4l7C�ABM�q]
H�F�N��깃Iv,�k84(��<�=�SHxq��#[D� =|E�a�L�jM�U��y�2\�������ժ���^����ht��x�U��j�� ���2��3X�=r�jDc9��|1\����Y���{2�ͯ`f����@h��S(hZPd��s�¸7��9�D��>ui��B��\0a@�P��Jo�����$3��P|}%�Ħi-�1$+2����)2�b`B7����0'�vzș��F��&�m�ÐۣR���#�#�x�Q�-����$>9�"��oE:�1͑g��{V��Ӂ�N�V����vXN�gov?�v�/k1X@�����gN�l����z~l�k.��Bk���0=�����t5*��?�pD�7����*C`bl�D#U�@���1��q^Tr >�'�#��9�V��|Fɠ�- �p���1A�7ds%�ɘ�O	g\�����qb�w�wO��@P�����$]ؙ�R�kK9����ԕ4^x#8J����n�xN��aV7��l�_N��B������ ��>����n��=��M�Vp6��Ù�#�G: ]*kC��]�Xc��R���an��#���r4d?��������̹{7�'ٺ�B��t���[u�İ�i�
BB����-@��BΆ����/�@�Y?N@��D�b���հu��ʞ����퍛5�w�#rm$�l���T��i�D���ih��z�����L~�懝q���ě<�I4�����,�k/�-�!�����D�*J���[rq[I#|v���PF^�d'��q�:��[��S���F��~�nd}�y���e
v�=w�~)/��l&R�J���#Uf�v�ܷ���
C9� �/t�
�?-��B_1U�Dw�?	��ZT�W�}�pR�Vz3��t�ՀC�5�/`G�)�?ʁ��'����[}�u�٣&&����pW�uI����md\��4���k�������/? �mH�Gs1}i-�L�X�Ʊ9^�J���-�c)Ƃ��c�.�;gڽ:�䦲��9�wrLBl��n����xW�@��L��S2�k��o��2�^	
/ފ��p@��t�]����VQl���X옓�� ��1�m?Q#�N[�������A�Y%\�Me�L�����y����Gc�{�C%��}[�	s��ʄ��^����P�w�Dh��Pc��p�;�=�(F�@�W�k��9t�y���q��S���-	�f$�uw�bԀ�l#F(ԲӮ��7�y�h��*��P�?�!����m >_u
�8�Db�^��0�wVm8P}�u2-8H��V��0�	p��I�\+��*��ֽ�L���A��A���JE ��{ y�`������B�7o�2�_�ڈՖYd�1w{�d�k������8���=�=Nn��Z�n'�!)ܴ�z�^n�*��&��ɀ�ư�6�g�Q��,�K/�٭�"`%�l����b�G�n�CŨ�@����v\t���	��tP�H���.���ȃ����H�0���,W�������Ɓ�0�TDWu$b�Z�!�O��|���zj�K\�vݚ�r�(�x!�z=��L��ƙ��_���9�[7�n.�}Tk*!?DqmkI�#�{�Wu8��K���,e�x>S���@�с5щ^����0KQ��d
�Ɋv"/� A���e���jK���Ǆ߭�!q!��a&}��u��E�~��gި4-���N���KEj~LtlZ���Q���3U��w�<Y�f�:x���)v���畭yV�2��E�J,2��.�|� JD|d\��h�#��'Ŝ�֥�6��/8��X(�h��_�i�l��KO��"\d��@��ڰ�v�"?-��#�&`@'�0�:�1��})�.���b�}��9!�Z��;2��tբ�b���d:��;WK#�]�|0�2H�r�om�t51d��e��d�Mc���A�#IZP��3uX@��a7*���m�� ����������Ɨ�o��[m�����k�2Ũ3Q�NR�ҀS��T�a��Vg�)e�t�=�������c�-x��V�;��e~�TM+n+�oa��A'��P^�.�%���G��*��2r	��������7���������yò�]��<~6r���U�!�q�V��R�q�Ȗ�k���b{c��W$�
B8�k��^0}���m7�<U�/k���1��!�q�g�ZÍ�ב4�8z``qa�p�����ʹ[~���WN>�T=����^���4�c��r��yh�z�����<{��Ңd�rj�N��0J˼����<H�<��hR�g]��ӏ�`�koϟ۬���~�
�LMX��X|GЅs`S�����s��]���c;w6�E�*�\^�,�%�p��&�@+�,�łd�Ro��T���xZ ɮ��:fù�jx��q�fD��H%1�'����<�տ�4�?�Q��9f�K�@0Y�٪���J���Vse���i&�h^Ef���HA�T�)����aFT<��,����E��)���9�zר�$�tHpz�%�`e��������Aڙ$,�8�<X���9�r��X�	:�!�#���"T'k�G���{��N�¿�������Myn���t�b�쪩 �F�;��o�u(�P�?�����P�~h�{/Be����/s3T3/̡x�x��e��Wq�ә�|�x�-�f&��6�]}0�ߪ�>�w�U���W��x����d�Ց#NQ�m�q�OJ��՚��I�}	�4��6G�TWǿ��'�&�y`��4htzg�����U\���`0E����Y�������x�)�(';�a,��b���tS��K�T�r�0W��`*�{�a��X�l�oj~����������d�:�J�<���9�0@��a��"U��4LA���c�xMs��Bg���%�.c�v���8f��볂�MA�`:�:�#A3}>K9[k�B�zp�(�r�a����4i�/Z���� ����<�V�� j%��Su��W
�mg��?�~f&��X�q��?��#�3M��E������$�c�~���'�F���u�/Qpz�c5�rG�����x�4��y�\H�Tfv@(�o��/��걧M)��]�OV�/��x��̠Kb�����1:%p�y�H��o�
g���ёƑ83ڋ�֩��K��H�nS�3� ;W���,�uF��_2�yc�����ԃ:�y��ŋh6JYm^�iIy���w5�T�%����������j��V���i�\�����)�?M�Px��)�
�M^�l�Y������pV����jz� ����[�G����2,oTW�⾺��*	�}a�3Bo��� �0��U����ʜo�0���gڵ9_�����������)���PPU�"��Pi��;��b}'�oG��k���o/�2x�U)�u���q��^�G`��qT�E�&G��G��ݖ���8�_���.X���4i��Z����8�K��MC�ID�VV�x*CL?�٤��Sܾ������Q��#޵̓fE��\��*-��|2xD�6_Ox��G��Y<p�������-�sC�7�3*�$�Qؔl'Q����Ol�U,���� �-̸�ǟ��d$���^FL�w���1Q
R:'Τ�U*�5?�����,�BG�L��t��П�m�D� ���Q���!c�"3�'�&���ͪ+B>|��ϻD�A���~�1�)Sf�7]@Y�ZF�� �pt`4��ȍk�|�y��m���]6�9u�Z�N�a,Yp�o�zȮ�◗���W���a�=˺jjc*��ě�mY��El���w�`J����և�D���ޠ�%R<���,b$�������JK|����Z�z"]�V��|��uv��{��B4̚�N���k`��!��#����{���O7�6��?���,o�A��v}��S���2d�5ʦ�Ŕ�r,�+}���qa�-�Ư��-$�K�ʨ`�؋<�x�������}�����~�QpL�qB�ۆ%m��PҥLCʎM�����X������FZ�T��{ONn5�k�?��f��K!ȬqdXX궩����&=� �N�����,��x�zN����zK$�!>R�i_/"M@�kғqDDk�J�	;�������V��7�/��vyz��\�\#�
Y��h��O1�'�\�'��覒;��!y���`����C�H7�	n�5!�9&�E�cՌk���-x2="ɮ�,�� ����}����<�L�k�Y�{m�),�= �ܱ�QW6�L������mV�b��K��Q0i:�#b.�W����96�����K+�-���ξ���[�����s�.��Ͳ��d����)��4't�q(k�/��/��f>�nikcZ;K׵��(�cs�9mQ�b����ӗ�/-{L��W�9I�T�܄�ڪ
_0(��N��Y��$|��l���v�9�6o)~}e)���警�BU�۶��	T���H9����%�~�ޙ"f���n�ȝ�Lԧ����`U|jXusl��6��z9���d���O�ME.?Հ���{3xR��%�j�t�o:�YF�Ű�@��Ї5�vg������] {�z�{JAW7���\c�^4[����l�Q�qj9��͆x��}���}����fֿ����a�S�ƒi�ီr<)��.��l<h]�{���8��"v�����KüH~Pw"X(Qv8��>�+ �����FDa�m�O�0K�š:cT㖰��T^a�/��1�EP�ms�g#�e&o��Y����:ʶ�����������������!X1K�/S��6�y�����x��&g曜ڪ��_h�������%	��$�Ê��^�(���HLj0��%���{Q��q�R���G�����π��lT��&'|n�ѓz�Y�ɞ�SN1�䧘�BMG_��ٸ�'��F���H�#�0��*\�`H��+��y��as�\B�� ���]}F���뙵끜�/:ZU^�����5�L�r��cb.yg��ԋ~������
Q5a9i J��n,:���㝊�%nx�[>�������jIh"�J�z����H<d��o!�g�
KЌ��_�d�%���7yr!�y�V#�ԇ�Q��%�6J%\FC��޼Le�T�c��|$��V1^\�k,	��HCG�p-��=�'��\��b��#>T��$�ųr?������}�21�%o5=����E-�+IoV�#�}�����fO]-{,�u��D��odl¯݄a~o�#�l�(IFh�����; ��ERs�~S�A�.oKE�Ȼgߥtf���	�Ũ��~��i{&a��G�� נ����4w6����	��g[�2�S[�7l��-
�%[KG��ȃ�T��jY$��~�m�J �r���@��NZT�4Gې� �Kw]�ν����InR8��7�	�NE~cB�P��� 	�h�༉�~}t���!��#3B�<p�D�h{���F�RO�ۏ��g��
����c$K�ݺT�կ�@+�I��?�������<| ��R݆�����L�Cl�5p
�sK�t�+�Ĕ�ʩj���,Ls����
P�96�0/ ��Δ�1G=ı�of�MY�[^וk��/ �e�׋{zf��:�<�W�8�8�h�M�����W~{�p���%�d��\�#�����"�8�U��t@�	|�Y�.'����yN����1Bu���R��Ŵft�1^R+��f�7�Yn���X�E#2	��YL���LN��K;�ş���4�";U�g� �IK!)ZA0��tvg���p�I8(�` {S�?80� �#k�vIW�)pm�0K�&XJg��e��*/��$�!�i�����(EW':a�\���͔�G"	!��2^j ������,��ֱ�6�R+��A(�[<��b�Ь)������19�@|�Cĩ$��s���,?���[�O�𺀄��TB�\�.�e�Ce��k':fs,�'�2u��/w}��;M��U��EJp�G(-� >�s�]���/���eaj���X̎!�=�u�����6�g�?��K=��?���>���hƄ��_}
-~,��,��w�L2	�S2�D��oB����x�?%J��'#�����Gs���;r"�u~���A�Ʊ=���g-�Ȃgae���8R����a���>g�Q~w�34[u�� ��Wғ5�o�^�����h����7k>;)4b(�[{J��	�qǢ�D�82��>���{b.`�1�3c�JH�
Bn�j�-Im���'������06��˖���&!�xF��pV��[�sG��M@#��B�6�þ?Y��T8~e�n��t\��GWt�#
�LB��Qd�܌�a�K9��sN�"���`�s!�-�AW���k���ə�Whk��@��~�[�ɷ]K eG1��R���f{W&��5@��MD���?�,h9����S>�p��CC�B���~%y�n�Y��uL��\��Ey�ʄ�B>7F�z�+�w�*�Y�-��͇�(yx$s���1Ӷ7W�B
nAF/��!��պ���t�bT�A-ɴ���?�e	�[��\w�r���\"h//S��"�,��d��Mqa4�\(�=!��g�S�ZI�E���*���T@&���H��:MB'�6N�8蘶�<���A,`���x;�����!������'޻�e�G;Σ��a�b�E�(uT�E����`�l�ZL��(M�*�S�f�-�V��a�#t�&�3ܗ�Sԥu��jm�G��$�h|�۸u�[A�ڃ�1�.�s��p�(tσy�)� oY.rH�����sS	
k9�t[~�]ۙ������	-�D]�A�K9�il�&*F~�ݙ�P�f�q�r���׏����[���	'�Acω�9�'(���ud�KPҸ�ME��G�oI��3Z����S�}�x��Ym��	O�3Q�c�Y-�сi�#�((�������{|��=FB�'�[��3��K��US(k������~� չ���R��LGK��hpB��5h�� K:̴��eI��<��Ԝ!�x;*/4/�('QN8�%A�U�3X���p8C�w�����Io��c�����)k�ħ�m��a���hLy)�y{F@V9%���8@]p��� ��ЌWJ����3g�Y
���c��LX,�ỗwR9���q=���l���ldɶ��ҭ7��������@�4�Um,_E�v�Uq$ �����H�m�F�U՝ѓ�g��:�6j�u	�6Cκz�!B��; #�6	��ۏUf�������i�1; �z�W�|�@�N'���.YȌ��+vY��+<̖�B��o~�'���(�x��\�k�\g@��us 9�������}�وF�Ǉ���!K�Ƶ�#xￇ��A���� %Ә~��R:sH����<�#�M�T*�=�%��Jt�����Q��=���}��Fr%��=�`�
F��b�9�ݎ4��miVޒ�^efQg��
��>}AT���Mζ����й��1'0bQؘlP>A�ǫ�P�g��}ϡ�Ss��&*��6n\�"z���2��dp�m�v���^|�V��PA�r�˿�>/)��\;�O�a'nXe�ЖBKo?��h#T���E�ځ̥7��5�����q�x��!��7��2H���n)#�F�j��	�VQV��3n�{[�brգd�x��&����?� ӌ�ؘ�>�CQ�>:y����%�C�uWv�P�vZ9Fψиr9�ds�E#e��߶x4�Z�[�D$�*�{,.�ɐ:�KP�$��j�[$]`A�u<�Y��z]ۊA☵��6�9�԰��B���r��
Y)J5-
�K��F��N�����c\%vC*r�0¦���YM'I�绾͆�\ hM�)�Ev���y�/:��|7�������KN�a�4�ךo�F�2�b �+`�86��ݸ�Ȭ<�^��Dt~l�FiB�j�+�ȫZV�"���F�T�(���\JS�u���V@z\�^���Pџ�7J�On&ݜ���!�	w���U�����MɃ^��X��Y?E*-�%����K�@G;�ǉ�ɣ���!!����<_�s��HJ���e1��p[P�p �-��i�^�\}�yc4��\|rE����zT���p����(��&o�[�P���y��e���!_����.��c�ܛ�ΩI�x�ʏԃ�^��N�4�é8��S��*ٮ�Ĝ��i�#��w�*��na&(��*�˫���2h�>��0ѷۃ7����	����	�lQ����6E���̢��Ij��u'��Lj�$9w��p���	����9�%c�c�z12�z��0Ȟ���v@������WFC=�J/�i7a1ݭu�BZ)"3Hݑ��UGY�3���N%P��^��@��"�kmJ�]Q\M����o&�x���sB�ۻ���~!�!�N�8\�AS�D���sj ;o5�p}040KUv��i%8�nN�ZG�<�{wt5���!�=3�ңQ?C=i��M��7!�#��dl.JD��)���C�@�/۱���Ѐ�V�_˺D�=���%F��p� Mx�=�o80x�<C����!�ݍ�gh�ttwݩ>SѦl���W���T�2_55�r*�ךRw%��Y.��ُf/s�����V�6�cK�6��мrE)����Z�<<,)j'�C�B��bu��D�㴱f�)���Z��o�l	����~��h�HS�\�>W� 6 1伱۔�5є�K7䧄k/�����n��	|�����p���x�D��lF�DZ_My�2eO\�/o#Ƿ"�B�M[z��]����D�������qA�^�5�d��@�%5��,���A���yM�-1�iMWkz��D*AlM����YD�̼z�F�����1p��Sv�Y&гr�沮o��4�v��4Y�nɺ�,��{V/�'9�(񼯹�����>{/�M��|�/��Jɝ)�8������k��i�M[��W����N*�-(�����-������M�ސ����`d���=��v��X�l��J{W�C4���6���������~��Jr�}>l�>u�G���,>�֡˶>!^T�:�y!Jڑ��UM,�����a��>/���o�y?���G	
'���y��@noD���if
l�qn�~���A�*���]|y�ͬL��ױ�#/l~���Z�K��=�2q�*�kzUW�'�������Ho�凙v�eM$��`f6���VC� ��:l�.v�R��[�S^����[�����f�"��$M��Vw5�m���9��3{�g�{l�9`-\���Z�?A�􍍩���!��$/�`���ͩ˦���������gu��y���<7�ς�>��J	Q�~�%�A�6�ٖ`h���)"h�2Ǯ��Leq����:	mM�n�\]+"�0 @+=�Vy-Xg��3�`��7�LRZl���X3*�G��gǇ�>&�D'k�>��^��kFʟ��)O�S/�~� ���d�
D�RR	�7,wʩ�&Y�Z�2�>j�x<�f�/g:$̃�YS0�J<7��D�x+����=�b1�[�.��LG׮C;�
����r��2}����W߇7o��7Q��2��ZO�����-1�gGo5g"-��:�s����U����V�;�86�`��O�+o�L#v<���A�t2����I�2H�M���@{Ǻz�y��L�* �np�����5��3Lo0DK(;��;��m�A6 �Nr��"6kF�p�-�� O޶���]=�[Cv��Ċ�� ��a���QS��y/mG��M�� ��Z���A���
��XV����∔6\���t~�2��������7M.d����>L3�ZIڪ�:o)���UueL#Rp�I��_��-�	s�)�*�B��7.���b��	VE��3���G;ұ!�}�w���$�֪q.�g��BD��ͳnp.~a���qE���Py=���ǿ	,vS,,=�/!���bI�-�G�[�<F,�I�%v�>'A��ќ+G�^���:7�T$�3�� 
����(�w���6�X:Ms�� ������PI���T�L�E����5�H����46�Ϳ��<߂�B=�5�Yt�ޓ#�0�$s)B:V;�"��bfE� ���y�є?G3=(0���&L�O�o���ܖ��o&ĉ-m:o��V�����T��-�6��7�§��}���IvX��7ƣF[WT�v
+��؆�e�������!���V���Y��@�b��_d���9��q-������l�}�ŵr�ٴ^Zw��=N�1��+[�}x԰��Nۀ@�x�R����xݵAF�~&	��gR?{�^�J�ZO3���$vmv���5;y�XQ�!���u"1�(�'����q_����ΰr���Ț���%Ҿ���&,l��l;)�t�����R>���-��^� d/�{�N���dc�;�x�+��q߮�h-�;|�b{�8�
�����ufML��=��K�U@I�5U���*���A�/����1�e��
�0�驲8���(Pq��k�z�?Q��f��.�E�z��6r��ȏ��!n��L�+��9�q}������;�oKq�C��&3f�8��AbDF��&;2���׶.��������Q�5Q�%s�$���ɳ��_�����PL����dHǧ36�tL�d̹Q�+2�g"W���Ϋ�\��VBi����HM�q�ףξn+áS�l�~�C��(�zC���e@t�N�N�!��i�yӹ�b�KN�|"�HX����R�+ͼ�k�:%��`݂��a�����e�%i���)3��\�:��KAZ���d<6&R�Jf�FP{�\�Ա"�9cr��3a����  N۴��u��f�s�M��wZCV����9�>����.��@aȰ"SAd)y0��̬8�k�xԺ���n����ֹFS�PY���D	s��е��%�����y�C��B�>#�E|�P�Vy���>�t1�rC��/W5A�=?ߖe��8�Q,i��p��9�n�+��:��L�O6B�_�aoQ���Z)�σ��j9�%xW�������k�<r{�6
ƕ�F4� B��G;�P����*O�h��B�$ff��ܲ,�c�0��w�\Nlu�i��p�g.�����;@��Ć��Pڤ+)WN��m�vד��Y2aW�,4���BK����5��;f8lrNX�9�&_�e���>�ԭ;�?�)�^�"�dTg����ܦ'S���W]�Z�^����?�$_{g�9u�Q�I@��r�2�� �`O����
C;wz2�Q��v���K����c��?���4ȽeY�+�����y�\��!O��O�Uc!p����fT���;dx>)����	��Qv.1�[�z��d}'����Rsa�M��w�9��.��&�ֶ�c�� $'�6��������kT4	J˘7R��T���yy�9Q�mx��L6~:���+�r����U@ݳQ�+SA��櫍4�}��F��UB-��9���\l�UA�;��0���QP�d��zܸ�,o��
1�qgW�!(��FH����-o�I�e�}�bݾ,5@�"د3D�9��z����fO��ꥆ(�"��с  �K��PN�*��lS�+�bg�S���式=�r!�.6�ӝr��44 9'��.��~���^�b7��������#?o��V���"r������RMk��?�K���c}{3j����-�r:�p�q�e��l�յs�h���Z�jE��� lp�b�`>�}*�P�5�����s��ǟ�=�����DX�y�:Ȓ��^�{�8s����U�=�fk�n��|����SL~�'5��H �py+�]rn��i.�^��ݓ���l���NXDoA�¼���wU?� �+Ǣ��^�'����]�m�Z�^&��M\���6j<����#��"H���M^��0��3jPخ��ҙ����u��� 8�Uk;^U�8�	�i=T����E��8:���?��ӟ���ua�R4C������I�K)�j��_hq��.�q��B�~�5����N$��\tC��TKCƹ�at�?�����bPw�ָݷTT#.�\��U�!�KO�m����'K;�	�����?\K���f�ӧ�#+��:���,7ɑ����P��e�B��\E�bF��^8xYe27��o4@@�0�i��p�������P�"���P}�S��|�$�Y*�]G
�n�����K��jǨ��s�ꞿ���������aٽ�H`�4����|�,��NC��g%:�@�����jG?�U;X'��g�S��#�A _�������K�~�l�!H����d,�S/<�EL[��UQUR������H򂂧1�o��N��E]{��ģ�9��.��c8�^93��-�TY��bڿ�U��1"�Jq�3r��/|���]̀�R��X"����6�k2�/����zV`���O�ұ�#K�j���߅:�c$���j�QǕa(/1m�Q���r�v���.#�p�3H��I�/�tD�ڤ/�ؖz+��c����D����9��^��eb�>�d��3i��Px>qQV�#�(���65�{�$LM�Z4�C6��گw���������Í�`C�[Щ��0�Z��;S�Y�����F�rz��3�lP�܎�.CF�⇰Z$o�ks�:^K�Kk��%)��v=[f�N�L�Z��\P�9�BR����Nn��f�Nt�����9���mV��p�Rƿ�2�Lb=��_�i<�X؀���Z�H��ԜA���mO�O�F�*a�<F��<�f���^��v�ۙ� �6��Wc�#���ePc od���� �j�Z6��tO�~y!L�АGN4D׆|��	sw�3+L^)�g[��1'��|{(Y�u��Q�Q���cH�Bw��8�C�w���+�R�F���teK�k[���\\����-e!�M\�-b/�N��{tɂ�s�nb�|���C� �0�2ښ~��2;���X�`�l�4��x�-���>z!�mZz�P�ę!�#va���(��O��	�sU�T-��&
8�2�R���v�Yb��V��x�Qx�X[��WM��Vht���8<�y0`չ7n "�7fB(�߉��D~$�'�8wEd�@��I3E������2 X<���������[�\R����U�̝��x>����e��j�?���&j��hW�A�G6gO���3�/�ַ��.k�ѡ�o���*�`�z�N���t�[����F8�|�xG��B�s��ӱ���"���3�aZڝ�����>m��|�I�DJ^s�O�E��[yL���:�+�1�����A�aЛh��:��͔���.Y{��Z��`$���8(�����vh(K�΄�_M�E� �-t���:������ffRC6~e���C�m���Չ�hV�ǔ���]�^N��Z;<�����:�i-�T=Η�C���%%#7�:�!����^!��Wu1`7 &��,o�|6;�ᬠ�ϸ�w�j���#��,�ۿ���T����<O�?��x �h����l@
*Ğ�}���FJ���ꎯ�dpqP��#�c�EpT��e^�
p�ri2��!��d�{T8b��E �H����A^� {�[�������.|��ϲ����S�;D�u,�C4P���u�\�Lm�*��59� >o�!cX��I����F�Smy0��t�=fң�eJh�ko=���{�XG���e�!�?�L	�����69U��~G�����:���`(?���z�t�7�:��v0��N��d c�
vD`sT�.5�6
��xV�a�_�+��U�UYJ7�+X߬�U��둊�*i�
��2���w��]���|���
���4��˨�+�e_F�w��y5^����i��Ɓ#�QD[N� m�e��՞o`�{G	��_�7�9���׈�����l��q//�_Wu���S|����(DJv�[l h�˜J$�*�(��u����4=\�D�k:K��\_Z�XTZ ���v�S�m�@[�͓%�P�.x��ig)I�����h�������ǱH������Ѹ�Zް.4o��S��U�Y�H�B"+�| 5k�߷���Li�����s���bB�n���p�'�-�SOs����;j�+�R���2_�aޮ�0l
���Ū?�|
a(�2�Dea'�*q,@i�Ao��\�2�;4�� �aPDKx�wh�|D���P_�N8]�-�En����F��p8x�~�ǘ�U&��o����6ae<���3:���>ٺHl��'|�~'�YJ��!@F������*�5�Ĥ�&x�M�2����E�iK��oj��Q���82�m����p��d�3�_�ɞ����a�V�)��Z��� ͨ�;���CB�(�����S^���~N���x�.��A����T����x���rs������m���u�M�� �V�[�,�"�[�.�-�ɨ�Ge�u�Dt6U	 ~�
M�:� �w�w�Ş[~�b���\�Je��fM��6:�F �q�;g�sr�w�O"���ң�Mq(���Ԋ�'"�?_-�c�טZZ�t��[��`1��zg>&��̈́"�T�|"��p�����y���ò��ß�J\����R�95v��;f��c'�Z�I=P�/K,�� �<1&VHo�J�W�S$WR�&󽙎�}iʥp\�2���9�Ł�Hq�;�
���_Y�#a�� �F\k���~٧�P�d!��5�q�������l��e��{՗�4�C�@j\;� X�����\IzX�� � :�LGOP��S�C	;{T�w�[�;7h�4�cb�&��.��jV�E���b�V�;�ϣ�sa 77{�d�;4:���L��'���	�:�����tBI��>�ɰsk~hE�m�����"jF��^k�Y��|<��~}�M��ύC¾�� eEU��U���X�W�Z�5+��CIS�Ke�cN���L�hO�a��s#��
-���$��}O���ko+�3��!��ý�}�
�/SA�г�$ʢ��G��P ����_~�|�������0�����IA��`���m#T��|"h*�� �W���7�����k����'����-�l��?e:��muˡW�ףE�T8/3���*�Jw9�$�����y����Ɗ/��\��m�E�@���E�/ԹЙ�	�	椔u9Z�<�Z�I�D��@���d.��c��R2dL�fdd��a"��(�Z=���|mQ�yO��f�B���%�;�<ea�(^�0ƣ3�>�&7h	���v���3Q>���4���l����f�먈a����zǶ�|�jU%j��nE�r
g�Č�b0�n����6�ͺ[�I�1AE-`��U�pQ�ʌ��E��𒝎�}
/�={��'*����[^��;��evo� �}�/A�mX�=�Q(V,k
�-|�����3����pq�|rg�=�[��w��~����Vj���\�`"���bJ�B�rش� ԥ@��B� ���a'E���� �	օǴ<�%��c�5�꺈Q�tY�v�a�#AN|�Sj7�sy��"_�.!�I& �?�C�:���n�t����Θf�N5wH�B��J�{Fu���ȈZ�����n��K+��ۖ4Ynҵ��=����f�ݴه�N��k��&���-%:�2�[ua7�Q���P������
�E���ڑ�=Vo�;�,P?���"��"F(-8�f}K�x�m���7ʮ�ݫ��n 1:^�sQ[���f����1��{Nx+.s1�o޻�,��4�e�#��< $��$��pt�6A�5#6�j�L](��Mf�O���T@n�q�g��L��V��[^SX�*�K:�m���l�w�P�Iz�R��sJr&�Zy�2��q^�֥�i�ԕ�Հ+:�]���1����tc���A ƀ>���85�0�7�ެG��J���0�F��'��o���=亇��h�j�ł-�;�ݨ�%�u-�ox>>�4~nƫ�5��k2z݀�Ǹd�|�QE�AEW�n�F���p*����A��H��)F��xb��H�cg���'�V�� �p��4?�8���	ʽ�S�@��E�����õ�=D��H�5C�~���L�`�ʀ�
�P�@a�ۯK�Q��"��*�2)��������\�'�H컙	k(�����~i/Q|��%i�,>%�*P6w�$���z�N���m�H�1Xz^�a�%}qo,K=�������̟5苔�v�S�6�&�����H���ְ�}�������ј�>�P�a
�hXC������h�`�&*�ɻ� ͟c�4Pl�|+.f��f�e��u@���~K�?�{R0��4�g	N��a�h�����+ЉtəK�%=�����̿b�j��p6�oc0���O]�I�_�z �ڡ���W�O�4(��&�EYb�ׅ�5Q>����������}�5e�@~��X�ۙ�E����@�:�C�B��́�e$�_��oY2�gaG�,�Y˘�[�rRN�Zh֠ʃ	Xc���;�-�c`Cuܔ�ּ�!WJ��R�EU="�go�,
�_@x�sX��a�X����1��c�[���0��ha8�D�b�wh���G����j�Z�Bi�s,%us+Kl��.����|JyGS�q~���y���`F`�ۄ8c%m��;%�hc�s?�>�4K�B�wXt9u��:�+��_!�|D�2��;����[��n��ָuy�Bk����,|�>�b�+�����vP��F��C)^�����	�'�g�M�#�?˿����V_�{Rΰ��5�vfVcU���O��%��
��� �@W��,D��V��Z5������{�C{"pI 肮��ݥ �M�'�Vׯ�W�`򇕢ʀ�$Ok�Y�|�)�����Mx��~Klo��v���}t�a�҄�38gB 4]�@F��i5��)8�� �C�����Ob4؄q�!C���M'���B�(�Ɩcm������X ��>f-N�n�V)���$$���<JE
N��>K]���˯+gLmt��`��v���h��d��<c���8ц���\��t9�8R��Q�}�L��eIgЎnI�]�J�Q|I��^vsD�����w����)5���1|kP�0O�<0M5b9!���:{tt6��V�U*���r�k�n����ϫoW{5��V�Z>RC#�h� ֑����օ�9��e�Cv�\>W�I�Y�
6������]��4B��y��#.C�C���*L:g�ż�.�|�S�L�����=�����'9`�t��&߸�;Z�7S Sc�rLL�fei������[T��8�a���(��y�'a�Y���#�v���V�_�DP	ZTDUU��,;���up&Y��% %��z����g��1�\�������s�`�خ�v��]�������2`�^����_B����6���E������/J ���NO� ��X�R�������@#�	0���^�V0{jW�G�S��tu4D%]K+e�#�L��;�q`^�xoT��è�lۏf�6pG�J���䶃�{��,���赻b���}�s�\�j](g[� "��8�|E�=�s+��YFI5�+a�NK�9��l�ğ���;K�JҁÍ�%҆���;��/F&o[�����w6_C"��W#�J^��G+���"u�O.�A�J�E�E�Af�=/���@��u���Rr�R=b(,�t'����7�e���*��l傭�0���#7�¼�v�uT���JG9g5�W%i�d����x��&��=�Hx77�]f��tJ�jY˓�,���(tI��ks�ҏ������j�GbN������7EKW`n��M.A�P�Se�RK��i�"!�R� f\?�ߤ-���@��B^�m�{�Ǎݭ����n,��
ä�K�TD�9f("�~�\�����U2��wB�E�Y�7�[n��8�D0��k�c)������Rǉ�z���G{���X�x5?�Mӻ�ܵ�&{����J �+�ۼ���"�ˏ��L��a�o�2�K�U�7� �ws0�v&�Cc�4�s�^��Tّ�d;�GcBi�D�Y�3���7#��LK+�&k�6�RU�[C@7� =4��҉�v�������&[��:�I9ws�+�#�!u]�"�(w��U�\~"�*/L_�̿ه�o��rQqy�A��v<�\I���D6u��=dGY��.%o��Ӷa*�U-��qS[�mQ@��!=��e�:]�_�[���|L��[e�R�����S�+N��*xGL5�)2v)�\҅�1N�}��aO"����}�C���ǀ����#���:\�UH\Ltj}�.G��|��3%���c/p�T���	�ea�H";�^{C@}� ��iY�"�����Y���2�����{~ubqDU���c�,�a� Mʤ�8��5����ׁ�=�ҷ���x���ۼ$k?�bI�HU,w�v�8#n=�
��*?9�V]3�n��f�`�MK*$�̌� 2�y����O�CzmU9p9�����0��M��g������NP�h��gn���\-�'Q]4[��Y4��y�}��tU�r���i<BO q�$E��`��=[�7r�'��1w6Ĩ�?l�Z����{M64�됡%�RXV��o�tݙ/�ņm��F0sb!��#���;k�kb��vC�#G�7څ�� W'B����E����9��/&���wA�"�ϵT(�Zg<#$r�L��\[�}�N��w<7�8i��炞�P(���������I�-�2
�!}��7�oyO��E��2����8.`_`|�u���ϔmL�N�	����h��t7��M�q�撘q�v�ȥ��j�^�����p�,�|{��Hs�=�)aO�R��CCˋ��ǋ�[�F�q���7����uy�d�"G� �8�553��f��T��xQ4^�Ɛ=��a��;�$Ȓ)���*s��,�q���x9
�퇍�dqEvQ޹7# �F^�A�<q0V�X���՗�zV�b�)x.�!�O;�/D�4����,M�����Be,��2�pͪ�E����7�i��d�qG�����de�:7gfy�hRʝSkt�C�6��f��*p��)��g��ĉS�T|i-=d	���]*�$��3����6�����e��OyxR�FI��( ����{K��Y���^?�짱��]Z��M�����Z�-���d̈~��2�I�E!�J{A:�! ��wMẆ�#��E_�h��-͎�1D�2��ځ�����m��Ra����E�iM��(�6i�7���[��6kj�Ʃ��J��x�_�ʧPz��dO1�(8{�0���I�����5g�Wt�Brz~����S�b�.Emi	!�A"N\��������a/��(G����'#��I���/�KHC�n"�:Z�S��}��AfS��B�󐹛��+�c��* ���;&r���]ڽZ�V\� ��F�]�H�$���`aO�^,qz���7���Ƕ��`M��� �����B9�l���K�ƺ�
~q�R�ӧ�he��N@Oc-|��S�4X��D��ۏ����j/��U����c!��3������3��(�.�7�B���ҏ=iH�(��3��num�0�	�q�*�\p���r���Y�w>�{�*�tU�+�&T��~���H�,ݸ؎r�/��u ��879<򡇥#]���B-�'A΂�}��k@��*��Hk�w������T>��u]��>�}ä��[E1��fl#Ņ��y�Qy��>u���ƕepw��³��}_QGQ��ٚ �]A���eOүqJ������Z����Tk�������1�����]���gi�� ���b�>�2%���k�З��,~�?4�\�+5댡
*��mM0s*	b�((_���&��>m��6�|���.�T��P����4g�3��<����;I�wAOԩJ��޲t��T'@\����'���I������nV��&��؟ ��Ѷ(��'���Uf�_�|bq�4v��T��zp��;�>+��¯��������Kn�v]�R�ɣ;�#}�VO�'�*�o�3
I<����p
f$�:KV7���tu��G�w�?��<]���|��p������bU>QE�|ȶƖ�Ф��U���rl��h|t�f��v��
#��C���3�<n�OJ��J�=���\�U�h�t_�Z.{\�˱��7�}/{�p̴�� ҳ�A�����L&��F�	d90R���F=������|cXW�(:\�pr�l4Þ�AZ}�@8�Oh�{�B�.�g8C����f��ID���~���^��3M���-U�w� �,�նL�1����;�Oq��_������v�䁙���������z��}�f����^���/�SS��i7A��I��M�}��� ��-x��Ȁ׭�j�ҵgM�[[[����b8y�D�)�<��rw��� ������/�:C;VS
q�1���ϴ�@�����J�ɨ�f
�-{*CV]�d9.K$3�����ʝ�PMT0���9�WE����� ��Q*���jm����m�A�����Ã|A��}��{7v�*vd�;�jF\�ٴ�F�}�I��Od���q�	ƛ�ˍ���~�YH�*�3�n�Ӑ �
K��nJto�r���Cp�$�ۥ��pf_WI]pI�<��[������h�G�ԫr�d�9tͿE��E0�׎wo_��\'���Mߒο�8�t�jti5���u�f�~?�Ie\�Φ���:$���a��@�77����-3[bC�3����������0��������>���U���QU��=�g�%�9�8	8�K>�5��.���H٤ݗ���^c%e�J4ςY��X\��7,*���MU ջ��+�Ji����H�f���N\�~(TQC�d�¾�پ��	����Ҷ�L���_�O+d�/�}�n
.��֭p�A184�S;2W��^S���,�Y�Vx����{	$�b���]M�9�e���QNە��n.ʥ����ToDZ�{������a�-���!e�L��{K��0�Q&�޲7�:H�5b��7֠+4�L@�������1zZ�5�ε*/��ŲY��=�������eX�{v����\^\���}��!�.�%��,w��z��u�G�Q
��z�%aR��(y�5�F�J��ހ���9��l3������_z]|g��|�S�r��2�Xd�~��̪,�H�f���H��	­}`gB���c�����������喖��o����*	���(ZA��	f���>`�t������Jsozv�yR��>��Ů�/]�z�
�Y2àH�A�<��l.�x"%���T,-�6����7�XS�Bl<n���tl��&�J�?�#�FeYPr�0����0�H��|��-O���$k�)z��3!S�U���<M�

��6����`^��Ρ�����cL&&��E�~2d+���b�e3v��>�7�?��|����'�+�^-�+�z�
���5�m#+r�p�N��^�2r]Q�~�&����T�{.�dͼTF�U���\2j|t�Oh�����\(2�+LQ���_B���M�����.Y+n�d*�D=�v-�}7�#�9u���)�c����C�Y�C��n
"P��(�K��O��ׂ�
��W�7�6�K�[}�j\�����n=�Pp(���ֶu���D����b�����G��=����䴊;�����_e3��*s�ZD��4y5��8�$H���\�>���-h˲W�t���ֹl,9�./�����]�2�,"�w.�x Y���֮����I�h��6���3Qh����J$k��c�m�m<�t����(��5	�Q���w�mo�\-Y:�|�eHy�Rn��ŦD���@��=P����;��s��_C�inp��}m74E���x1NJ�j��Q���Μ�6�^$΄N��I�|�o��%��Խ#mс�����������Z�;j�]���+�h�ͥk�:�<����W�8�(��
������t؞�������{��[}�W"�1XP-=P�uk+Z9Uk)u���=Tw�X�WW���B
wPƉ�W�´�W�1����;m>��<Y���o�R?"蚁�	��0X����%���A�+=n�MR����~HIzDN
��C�������CA��C�*N�^l29�$�i)~��G��?������
7ѵ��	���֘��,v�
�^`i�675���D�~��qkT�dL����̯f滦׭B��G�kZh�֑��B�<����ey@ے�I�<�I��-��~�)cD�W!Cp�Y|��@U��;j'S��J-C?�^�s�<Q��=ԁ��ɚ峗�´�]`�h���U�uF�@�NY���zԄzz0����FbzQ�����3J��ߍ�%�u�����\�si���^��M�{���'|߅��b��-�'�{Qڡ��DŇ�����S̉��[0����j�k�+��;:i� ӻ�c=���i�T���X-�BɆ_N���	o�&K4[h�e��%�����o�py������w�3��?k�m��̄(��Ԏ���KfO�T�}zdi�Z<�a��Z�*�������b�v�*��̈�>��jpiP	��b�v��g�#�]��E�:Mǚ�%�Ë��g�L_���M�O5Ӧ��y����q�;5��}�۴�7��J��P��Y֘-ؘ���&�.^�XE�Q�*(�Q��tF1��Z4)DuS�G۪�qWM��g�'�0f����V�2L@�i����nC���Y"��;��T�)V�]5V�y�t�r��q�Њ��2�za��O��HR���+Z`�K`��2��#H@������YyUP $5W�PA~lK���x�ܳ���U/�+H��q�m)7����3�y]H�^$Ԍ�|�ʃ7�{��PC��ERd���y�F��lR�d�*�e��ǀ�U�!��7�os];�sk��Ľ"$@6���F��>ڲ��w�����tz�Ҧ,k��)��<�>w���p���+K���Ch��� aU$hQ��#=�E�W��TA�L�)Z�G��T�T'O���3�+>���3�Uȸ�_@�\�P*��k� +���r"2�H��k,�F��Z�����F����iA�����R0ܱ��ɷ!���Y'��eg7�]�1�Ah,��$i�׻��P�g?)�P$;S�4�B���%K�ګZ�bc�SOfT�+�n�'7|�T#"����0Xi�.?\�E��m�9�����C���d2[���:W��·[ě'�*P��z����w�^_A�GM���^sdXX��N�5$H�*���|9�%3$M�꺡0�"wN6�Ύ���Ɋ����qËM҂��!��ʠ���/�8zC�?���]�&65T�)@�����}�l� �wPy�^���0�q���dYh�{�3�z�r<�=�m�_�UD�v����� ]��١(����+pvHjX'��88+����R���W$c���<8 3�Sw}%ݼ.�s=��/�<����� v��!��a^	<~���5Ȉw�R<��m��a�;��en��`��S��U
0��/#�8l '����Z=WZ=>���^��b��M,}�a:O�F��x�K�!Qk~�Qiu;)N1��/������~z֑��0�FG����צ��փ0��l3gݖ�S$��ٰۛ�T��6&�:>���hx�+��7zկ�#jc�p��?�hW>]Ts��,�ʾ��x�7^���v����$)�����u�	K�"�t�Gm�L�N��,A�ס5EŻx�0ZR��S(����c�ٝ�ĳ��,��<�!�^LLh�����y@p�������U�~����D��9��S��v'��O鲰�a�8�]��,����H��G�[���p�T=��m$Z�A:���[�V�)�>&�2&�=4�B��	���XI�x��`$2Η�=i��
(����`=T(^�:�x�}������:���Ǒ�8PJ��?���k���hs���[b��dA����I�^�S�ޅ��f����t���H 埕P�C��0�F])�Pd���VZ3��T���.|����>�i�Vo=�o
ѯk��d�X5j�}����@���*4G>X�2l�]��?߱1��C�Nt�� �佧��r��stMAU�w�B_�6�qt�ZÖ�d/��aG�r�hέ�,+����$e;�1�~L�=��-�(��+���"�M�v�?��O¨Q����u$���LNu��ʩ$.c��5?HR�C���g��g�d�a�?]c�!�;s�,��th���%Mh`�(��e}��U1�� o�CbE�"TVO�*F#l���IVè���ﶾd�i쉴���F�^4n��Cya��a�ǣ췊J��33�e�_#�-/Wq.��D�uS ��I�Amu��ӆDp"w1fx�H�$I���-o8�D�-L��K��y	�}�X��˅��T�޲IK�L��e��s�ʾXsj���OA�K�-�9��x<������܎0�CQ�N��� �i�#LXF|�o<�+��&GXq-�*�i�����0[�����+#��`9#h�*X��n$�y�cN
�{S�����0��7j��&�ׂ4��K��OY�a� ?Y\�8����\Ԅ�D{�A7j�n��§q��r(7���r�耯�3!#������Z�a��������|��5-�K�3�z`�Z�~��J��LՑ�bb8(�a�7�"y0RUz�A�dXL�>#� ��IJtf0���C|�c
_{�6%MSc���Ӿ$G4�M|<r@����d���ӣ(���Ư�|6�ub�ː��9��"��	�+�� e���*txD�w41��*���
SOjL]��T��3�e��j��9��Qh�ذ-���9�g�l���Ť��~l���S��ނأ�.�Z�����m���f��f.Ƀ-�?�S��>i�w"F����l����Sl�Gi�0����e�y���`d�p��gW��Jl�W6�8f�S�������M�UY�Yz�p�@Z��F�^b�FΉ=�q R�6Di����w/������{��B������ť0u:dq�9w��a�v��w&
��-�8x(i��Ө�����Ew-F#@��l;�J�ݫ(Ck���˦ܤ��ooƕZq�!_�����>7�D>߮�e��u�.ҕ-0�p�>ó�Yͧ�i��ڄ4��k����́��O�n^�*����G�[=1)�����'{�q����(zj|}����*�P��c���83�J �ŏ�|�[�ܱ��h 5%s�������B&���_*���ެ_�&��t�7���ً���g��.��h����\m1>��T~�N���//s4��r���d5
�c�@��1t��k˂>!�9IS����aJ��QJ�Ouy�a��+w��+���oH;���m-%�]|wȥ�A3�e�{Ψ�&f�<#�n!��(kkN���%�0E^�MO�# π��Nz�-���]�J�9z�=3ˮ��f����53b�6�^]-�@�y�Ǹ�d%)���XZ����;1���<t������#�]X�Caw��$�w�׵E����C�M2�I@��"j�ς]��r���b%hZy�z�b=6�vO�J�IG��'/�_�w���d��y�F���?z���_�h�Y춼�����T��)������kdӘ��lfmPB�>���!A��0x���PiQ�`��8(�X���p��g�R\*��"�MH�*�6��M�8���m�f�������cd����e��q�[3Vn$�%'��-"�+�B��7�?�=�B�7ZWO��3!��'������c%�^ʕ:�@��?��H���4��sw���H���tຆY����E��=v,�]�ۤԊք�Q��Q��O�EH��Z4��Q��L���
��� �u�����>��{F�'&MR�X.�7k�{�\̆Ɛ��{�ӏfޅ���>����,{VR��JQ�M'�+�y��,���Tm�);�Z�07��H����l�ʜLH��	�P��(�}��M����L�N��|I�xr���S):�2����xJ�=����p%B@J�V�3\�V�,�ť��5����bl:�V�|Ob9D��/lO��M!���EK��6��Yݙ@�����'c��H�/"ԝ���L*s^�#U�}v���v������;]:�9��=�&���Hj�5���	w�xB���5�Ɓ����.������)u8�;Om���9�s��t�E6�׏?B�!�P�8�yqj�V�B����b+�R|D�\g�WXL>.��i��/������[�V�"x�w�;���\Bè���S�B�e"��)�=&��]�4�
T�M���ңf��O�:�M1BSg�,2��t��<�͎>"hy�DV��]�E��8��	�~�Y���u�A��Kv�[Z+(b"k��6��A�'�R�#r�>���%ON��FS���S�=��̬���J�[}�b4�i4~��0ОMt�xD��ơ����ڣ��{0
�	���u�##@��"�N���<NJ�4=����sF��4YO0U������Pquc�Oʺ�� �k�ЌmYu-+�7_mZŀ㸤���a�f�v:r&��n,HC��fν���/����� �<(D��^�}R>�ٱ��-�\�c8�����Vo=q����E�t�ŃH�C�g-uq�k#v��X��GMU��]ڋ�Qy����M�ƇyIE"���X0�8�O�]u]�8{�\$ ֗��f����[Mz��@E��f��X�I?��}mz�Z��ZJ����)��E�ؤ�Vr�l���b�d�!�ݴ�|���-H���;3_К(�8��G�f�/[����᷌�F2܃r�ң��Ngy XC�O(���#OhH��
�����~>�6vj80�9x���Ŀ^�r�c�	��LeU@ɼa�U���8���l�������р�Ik��!��J�����)�%�V�Ͽ>e9J��b�:�w-q#���+�Q��#�I<Jl�N�"�ھ2�P��\g߷9h����A��Q�&�YmM �P���vR��Q�9[�;��)�Ѱ��#(�Q%Z�ޝ�R�~c[��|A�o���`����3}����*`m-�ܪ�h6c�!]?�͛�Y)�i�=}��ԥ�nC���T�U��њ�g���c����YnyD9��FH�Ƿژ.�Z憁�\����%Lρ�jB ��$7c���������;�:�ht�܋��R�%��g�	J����<6xdE�	 j�-�� ��J�,(v�]��G	���y��������ƻ�k���×��~��0d-nG����:S��.��E�}��e�,�+<-�=I��}�WS6J_ޓ^;y��7.�Ep�����)�\t�˘c��f�ĮNrjٶ���1�Zz�\Ǔ?�^YPJ鼯���!�� �J��x��E��}���q�����`�<M]G{ ��ͦ�vP��7�����p0�N-�F�sj�:�Ws6����e��weFjJl��%	���R�*h8T����N���%J7X��v%=�>���&����g�Q���jΑ�J��#s@����K�����2�jx:�e"r[������;�K^6�.F��r \50do����J����"����NR��դ��/��Ix��%<,������w"&z����Ԓr-Q��s���a��Z���\�S�x+���w�	�ZNO�ʨx鿏���޺t����!� I���p�1�澅����s�Jtg={t���X�����i~)�_���E_DI��c\��}O�ۥ·s�yV'F�?��j�k5�Q��	=�ܑ�J��~Q�p�g=��]}t� �戴G!	!eF� ��͗�����;�MX`��?x[L�U�����d�JJ-��nt	�\O��'	W��blI8qP�/���!��8�Nn��ZaNA��9�m}�?d����U�I{1W�InP��oN@�_�t�X�+؍�c�=C��:����0�	�$��OfH�ӊ�"�'W����[�>��		�wj��b`{��z��Z�x�liE�3���rX�OU�z�|$~9�(eQ�&��4��7��τ�0ژ��nI,^�.��Ɯ@�0�y�*��,k�tD�ɒv����s���ӷ��FFdH�$��]����(�"_�"�o�%�?��4$��M���֘���rOd4�M�o+a(
�l�Ea�	��"8���8�㷯YB�([���K�F��JĄ���Q�Ɨ��9g[��	�j�Mr�I�K��S9��'�����y|�@z��zx�&�x=s��� V�e��m}����{Aey �꽁T(9�*�j��2�s:ѧLTj��񷣌�3�_��V�f/�H���Gg����>S���%g��z%!'p;_����?�dG P	n�����.,���#�3]&Ň���FB�[/gE����R��`Ҥ�8��޸�s׮�9I��n%������'�!i`BU�@Q�!�Ġ�����1���u�5ՆB/ʏ�ɔ-1��l��a���u'��;ѯ�:����7'�*�Zw���P�4/J%!�eH���3�՗�<���ҷ����e�@.�;S�+�"��7���Jj�Xj�� ^%X���5>������0I�����٠�ܵ��M��Ƀ"����P�|������?�����1
 N��cye�v���܎��b�eJ�j]�Z��F���vL�f_ˬ7�i�s�y��,��W`)�������)=ϧ�7��6�
e���Iu��8����ەlX=�dk	n@�$㮍��?�o�W26u�U������4�$Wa1�&�|?]nN��i.ô�\��|,͟zDʪ��A�s�Q�"U���gj�q[�ZP��O�|�@��xllo�D�;Zݒ/�4�vS�.`"�=
��wd�#?���#�<��$}>��Q���?��%H������������,8
Lԧ��6�S��G������q:]���m	�ڻ���{_��Rgs���̺K#��Q�����n��m�.=��+�v��^E闰?((�����{#�*�^��͘Y]��as._-yZ�K}x>p�Y�1�4+ֽ�2�����*xf���f$��v��ͣ��ִ���r�9����7�c��,^��k�߮�p�wϽk	��ZkoA�<����I�c����J�4��Y���������6Mpm6��!�+:pk�s=p�|�vS��겋��c����N*q|��c�