��/  �d>$Lw�e�,]�b�sᗸ@[����h/m<�=O�����M�XX�+�*�Ͷ�����,��8K��I�Z�oL�q̂zC���"��ǧp=&:�ZLW 
�!D�y��_�fM&�L��_������$i�Uf�@d(v���Tc����Xr�][hP2zTa��h����!I�CR��c(^�!�~W����B����Y��g��A�y[3Ղ�㲕�������ч�/tsn3������G"�bb��fu2%P ��ڹh:�~9CG��ߤ������H,��!әj�q�
5-����g`Hv���Q�<�ZR��v�����C@kl��~1>"i��b�aް��X��9U���-�ÿ�GO/1��*��04j�vQDU�J�����B�₨>��q�5,�O>��L�֡�<��P<Å 2<uwY����Ğ�O�C���-Li��bRԡ�r���ƨ�"��4�V*m[���D�+�K����4��MB�@Q�J}��P��5�tG����h�ݟv�/&�(d=�+o_@ ���U��$M��2��:E��պ2�꯷p��\�sD�bWY����	*��s��9��u�,�L��w��N���j�~�v�N׺�,E�V�[cCR&>k���dh��WQx����ǎ	���`xW�
���g��g�}�|%�f���ҙ[�C�a*kk�ѳ�n����	�
�9�J�
[>e���ӎ��*���t��ʶ������ΉsloBJn�K�tr(~ܯq�DOV3Ϳ�qߢ�k��@�H%"�
�$��U?��^�\k��eֹ:����0n�=}������f�I7?0�g^��K��L��p<B����D�'���*����M�{kH>��)�i��54��("e�;U�J�Hc/~M>��@���f k̎��)�Pl� K�}�D=�%�p:��o2�������>� �[a�=�^0���حgM]�o۰��dj&G�4��#�`~b}ԣ�v^ ���Z(GЖ�7��z���U�#S��W������&'c҈6߶�5�(���k��y���z�&M+��t��j�U�����XvPY���T}E�?$eY\oY�s��Ds�q���l-Z���`�@��Eǭ}]�ȝ	�ʁ�s@�f�b�Q*�Ű���Ϙ�@��Aw��ŘR�	
r�!�A����/=8-���@=j��e���շ��xQA��h]��ة
|�hCU�w��;w�������+�؊
=V��(3V���S֮=�|MTmt���ś1?!��q_7���q��,LY��h���A����tM����R�`̉mP=�����f�.�DC��h�OFa��i���	f���@y�
���辅ʾ���j>��?3M.3��mO���G���S���D�I����w�P�~N�(v�����(K�bO&�A��~�����W�]����	Y���d��H�e�ޚ��[%� �\�R�r@�e�5������ደ8Z��狉��,㾍i?���RO<����e��b*q��G�ؑ<�'���vه�ع�;��J;WZ�s�Fż�d�?&�zI
�ѩW����=w��OKE&{@^���Gg�\��&�}�U[9q�6R�Ӎ���'���ZU�P��M	���x�$����g�Mq��I酡5������Nr��oI0��ʖ!�2�lɩ)L�&�m_n{sϿZ�ndt��5{W)�?�D���co�O��e�\'δc�=`��3uwep(��?	L�)�ւ-ʨ񊣯�l�U�A�_
T%	��X3'�!2���/7�U��*o�˄� �2��*�"=���E�]V��f�����DŨ�����}�g���E��U�_�6��@(3M}�C�h�.�o��vg���0 �Dt� c�t`{7�ִL'�V�WC���%���O��ɨi5��<�6���;o���+�#-S�̆h�C��З[�0Q��s�L��J��� �0M����Q���ж�fT��[q���y'�5�[����|E��Bȼ����!�.s>|��A|E�2p����~�����경�V1	��W���`.1~��{F��a!�c�O����&g3�?S�H�H�ڬ�{��B��\�ݒ�����2��[X�4-�d篸�����l����w���ÿ���d�쐸�L��w�A���C ����Ǔ>��G�i�XI'BQ#~�Éc,T��j�\����b��k&�!�B�ù�du�1�Q���XG#S�b�d���s	N�v�Z�������r���MI!���.��j)�A�uy�2����3�br��L�OA�,� ��"�X�!Y��'�����ITH�z��z*Z�3��j�R������{�Vf�p�N&l1�b+(�����1x��)3��K�-[������ɯ\��5�B����i��<1~o�����<���{���,']D;������^���*����"!���0!��,�.+���u2�R���J}�hAeJd?oa���x��&5��^3��+�����qL$��v�s�!�	��7WMcr쪆��}��T�-�'EHK��~�:����).��n`��*�k.�/�YcY�s
�zi'o5a�d���W�S\?ݲY��\����l��R��g�R����"M��9��]u�P�z��n��n�����x&��sE�7Wt�1�&���	����,�t����9��8|Mv, *�iS�Ҵ^��%6yb�J����:������Q�d���<x�trf���$�X����jE&]i��u��ABÄWGIW�p��w�"4�� ����*�f�dc�<D�?O����(kܸ�o�S�#>��(�y -ճ����B�Z������VԼrb ��`��a:��|ɋ(iǹ@A������~<�g(k�����D�3�D���s��U�Q��quȽ��C�12�(�Z�d��;��4}�]�n^��!m�cƝ=�C��4��0�-uz>9K�D�����>6�k�c���,z��}�M2�f��~PA���+	�����M�4m�.?(��N!��Q&y �����=���NLLD��TA*�l���0 �"8�5���i���U�^
KEc�X�9���s�m����2���ⵡ�e�E�o�A[���A>�a4Z��TJ�>m3A�pxq�%s��$�Ιw�Bl8h�FD�sJ
{�G�^	C�H���	.�HWc�� J�m��#���YR��C\̬��2��ʮ���W�D\�Lw��N"����P}_�����K���Pו������@����KN�4�G����̑�bO��e���\�5-��]�s�I��/p��HH/����툁�T0X!j�%�wӄ�\�^Ϻ��N���!軍xď.8$s��/]�d�N%�V~�ҡwr�+�ųM3p-*S+��K�9P���� @�(q�Gx��Ŝ��� �[��yaiXB�Z�?����A������q3�Ɔę�� +�mѥ�Psa��ׁ׫<Z;�"Q^�!��h9qV%F|��:�G� ŧ�5f�Mtb�%`D:#����5R
7B�������tes��2�ʓа�3\и�� \[~F٦�K18�cE��dp�� &��Y������Z����Y�d��x`7�~Ȥ\v���D{�@�P����iqk��\v�k�����E�d:�����~r=�G��\��?�XV���Ndv�Z�~e��-���^�x�ϑ|MyY)c�*~��d�=ӻdދv����N��ȋ�e�}%Rw%Jʒ.�F��iHhb�md�c���-�!t�"�U�\K.���j�#�G�Z��"�� �_t����8�G͉�;rk���ۢ���Ob�\p��߼.�9R���sKc�Ca�n	�2���p�b��u�ߑ��$�.�����#��{�&���;���x*=2���>��+�������o�1	YR!�������D�s��:���c���������L��[p����l���~N�ty��뇺I��������ZA	{�ޔ�E��'��Ē=�r��`�m����v�M4�!N]��T�=S"�R�K'��
k�\]M��8��e�/���%䗶a�d���Hg��4�䠟���É'@� �)m��b��H	�q������]Rp=�1�x��,Կ!�dɎ|�
�[�EM����U&��g����ؖ0��;���#��i�l�S���S�>�{Au��L�9�螈w��i�>��J��c���i��L�W!)%)�ǋ�`	�ogU>(,i�wL�������$w�m5��9��=�*t��C���6PNCmF�R_�e���&�N��Ҫ���]�i��m3�1��@4����/�Nq֥ܛ��)BG�k7R/�'���5�>�V���I��b���j�Ц��OӬ��fvM.�gQ@�RB;^��.#p��'2	2��Io��RD�<�� ��̋�~�Gm��Y��>"mȝu��kuYTV���6�l뺞i���0Q͙��}@����<͏1/�n~�j�+��]��}jF��;-~����%������8K�H�~�Xuq;�'
��'\�`�i&�?��&V(�d嚄e��߃nF�ƞe�·�%E�������u��ZU��ǬPl�� v�@=#}��Pu��5K|	��i|oy�YF��+a�^�q��O��B�N�b���j:0�	Vs���=�^) ��M��?���*s��E)	Gr7
���dr��Kc���N��w��;i!6�������M�@�Z	�0a���J|�
��:7X���kfR�Qε�~�۱�E�&F���rR,���KmQ��,ȗ&�|�j�',���(V���}�Yεj�$�#@��D��V����,�	k{����̥:ʤ;��.��B�Z���ص��)�E��*:u��`v�r
n-O�3w���S�x�BWw6+p��!�����c,�
�c�a޴��>p 7QVdq�s�����>8�� �U]'��a��زB��x���^�n���C�̜�`@�;�J��1�"�XT�N���	0�Q^��׹r
���ok�Wi�l�f��s����ꭁ�I�Tu���y����L30�Ruy9�,�8�0���^J}�JK�2'kU�+��ޞ���L9��K��F+]�h�S�|�Ds1ǾzY�@Ak-sA�@�0�9.5i�_�3�鮪��!��䭽�X��4:@^2�7Xr=W
��b�*���;�̻��(>JOp�-�w�uv�ƷpYn5��>OH�,+F%}��}�� p�*���qz��V��8I���ݘ:�a����!(:<S��'@}t˚,�FW�e���h��*����w}�+���	d,k2�����i�(�g�G+J'�aV��Ngт�h�^�q�٠��C�
Z��^��v�$LV{��Σg)�
n����sN��j�N���D
b-7W8��#4ӂ�� ��s%�FQ��OF/�W=�󱎽c�5xn]G�ǳP��bC6쇘��0�w�s�Dx-��RI1:*��Y1�h�7�A�}�M����#s����Ϫ��GŇ+r��h����	½���H�%ݑ��x?�}*���_�7Ga��>1jLj@��S��C*��v�zF�b��9�fr�L�BH��a��aPq,��aH{i%��N�x,��܉@���8_����T�a��+U�SF�c|�.�A��`e��^k镇���J�!fd���,������=9�AN�6a-!�_(Z�QB���[�,�T���g~��G,��G���Ef�JH��I�-�K'=��8<I#��ɑ�m7�e��A�%&~|���Q�7tJ]����x�������(���R�U;[JY�N�":�Z�����|�5Uf5l��shZ����+��vb�ND�N ���V��f����
W�{8U��C�3ad�������sE�{��5E6\<=z_ ��	�g���Liv%��(�>%H66`�)ȴ<�?���[� ����]�y�Y����Ea�r�hX�ч\k�,8h^�9k��禟��"P��S&��;�o���d�@:����cF]r���4���iM��cg�����Llh��[G��}OC���X�O7�!�Ѓ�9`s
��?� �~��M;A���X�� �E#�c�gLn��l㈁킸���bW__91O���k��㫢���F�3�u���E�:�*�ڡnW¡HQ�7W1�e���3��{B��:�%��|��z1�I����ƃ��}��su��GuTi��7Ö�Xn:a�(���~���<RUZfUZU��F�����uhU�`�^��
����Seg�lMOCB�����$H��6\u6��+d�H8����О]fٽO=۠�a|�r򓟯;��aZMX���b2>�l����Z[wâ���ύո���oZ�u�+*W�F^n��(� �w���u���U�w~����Ha�������Cz���}�?�R��F�g�w�Z�2�����f�n�Nu�>:�-t���ڙL��bIH�	��rJ�D�_��2�{������	C��O�>Һ4W���f�N�F�c�����h�&�k�+*�P�{�ɞ��6�L*,�7��p����L u�O$f��[|ݔ-��wn����НR�v*�mC 咦��?��6����[��� V��Z�H���犻H�r���;������a�����1�ӗT�0,W(��*�a01��*�~3�u��)ܙ�X�(�j�ގ�vП^�
�β�M����l�|*ƞ6�;��%__	���%���#��:6Ѕ�+H�yi�"+��� <�J��� M~�������!��a�X	�iٗb��-%d1�i��U�&z��<D��ƴ0}:�[�f2���^Έ�yAR�j׸;5��+���sC�ˢ�<�W�2֌ū����J�)����#�v�T��@��Ly\��EE#�R�ZB�[N̈����`}nG�@G���5F0e�o��;ű^�;�1��te�#r��3"����<h�B��a7��̗f͊ײ��A�c;?�#UE��
�R�u��[,Z�'g���!��C���ˀ��q��u�o����Uj��{B;\�P�*�tH��;R��^$)�/J��a�S7cں"K�,n���tq�T�K�\1I�G��&���71�N�G�x�kR�R��-��,u,Q�.A���M�b2�>�zt��?y�:�5ܧ���LF�C(����t-�/�_׻�:\!`�LTՒ�1��#��+��P�;�\�庛�>Ԣe�غ"��7!�f$7̢>���M�f��!IQ ǘZR%t���Ko���6O�U �`�1ղ��������V�Z�� ��%c{�!�i��7�EL����*����
�^�4�hH}j9Ϸ�/DQ9���/ԉJ�
�!�MA�/��>��?7�iw�G)<v�|7:OU۷�djԏ8a9�'�����Y�=�&�ۢ9�gK�`c��\h^�����X�t��.��Y= $q�T��(%��II�X�j~v���,1x��U��h	+� Y=���t�`� ��`K�?
PtWO�Θ�QJ�0 ��)	�T�]�$~��+���W�K�f�*`��4�/�X�J�#�<���1�y=�q�F��u2�o\�Ɠ�/w� �^�B�>������m, �\����#0�AT�W3���ׂ�0'�~�4?��"�;�!
�hZ�¢AwО�2q�D����֜��H�)/6��'�J��߹��K`���cq�&��iӬ<82k��Pk/���r��u��c�g�1`�{���B�:����r?v������"�e葕e��9�9���xٌ�H%K��:�v>;x��Wm��tT_�"G���m��ݏ�%X�u!E�fL�)3�IہJG��V�R��P�{�F��b6X�[>b.?/��̯��a���Z���w�`.�bk��m�|!��.�����&GU��+��/�k�Ҩ�s���ۖ��X���2Hs�W뗝}��+T��9u�G_��`�^�9�Va�[m�
-�gk���Š�
F%����f�]�V�Iʁz�g�.J����sH�8K���XwH3g.e��v",zs!E,)1��A�{GA ��[����,_�t�_s��r)rJ@����{�\ ��"}+r�Fw��ΝԢ0�§��m�w�˶���ⳣ�2ua�0�����Yн�e����b�wz�H6��sDt��S
��B�!DD��[��~�ek����61���U�V5��a���W�s;�aX�:�a.�ݿ�ݻ���*���U�L���f<dl9M�K��}8m�dKh�5� ��<KGCmh����)å�=e��9	���W@�~�6f����N7�-�`�[;��Č�b� �'h}wZ�\v�b�
6q9���c�s�K�@�;�B�N�s��,IRkK�������1�s�:��@��c8��9ˉ4h�g�cƃz��s/NI6���B<���� rR!� ����͢JC.�U�
�:�}6C�N,YRS�Ǥ�&����$��Ar;��@C<�!�d�,�L�[��
�I�ل��cmx����3���M.��Й����3r���-x&�:p�^l�2$�Ѥ��������\�U�2�%S[�k�.�N��v3Y�lQX�8z�_��s��/=��LޗzMCk�������FGWb�ǍJj�����Z<�2q��d��?UE����"�Џ�'�m�P1*�
u/g--:�D�r߈#a�.`91�'�o��#�Đ���S֨��u��A��FFxh�/���ʅ'�j����� �d�o�CڿAp�S�l�4�*��	�"�f���/�n��a�:�Sn����F/o�+!oo1%���:`N�{,��]��L�|�qJ�j�y�����` ��	4iNJ��1%I����K&�����Us�= �s:�f����<��iH/���&�8Z�#�>��{wC�peT����S��=�#����{�Z��˿���39)��Q�V�v�D�1��]�U9� �����;�g����[-����~~("oYA/�1���D���s���#�M)�AH���\�+�j��G��ݙM��O2�P.�Sb#K!VR� ���O�?:�t��~6��[�)#�p	NŅ�Ģ�V|a�p%�t���kB.�1(���aA��x4aPԪ7�5��(�5b�|���q�ǵ_���N+1��cd$Q[���D_��Vf�3
��uy@�s
X ���/��5Sё[���RO�ﵯ ��ײ�l���U��J�I���õ�
�&6s�|(|�Ȩ�����EZf�����g�5J�"�JK��H9��=�F;��aB����[N�t��NC{d�����j��>��������PP�ž��֩�6�PY�v���͈t��FS��%s�K6���~�.Q,����ZrW��3 ����ɛ��l��x3	lW���I�X��}s��+gl�Ī�5�ʥ�O�ݷ:�3u�J��rg_3q��ֱl���w��鶼�KX��k���E5�-��ܻ�N_F��`Dv�@�?�/@���E�㶒oY�t��RRå�s!�}�aS�nz�S�lm�Ѵ��!��PhE��Z��.I(�i����J�<�d�&��5�|B����J��u~Ê���I�m���ZR�K/�l	��r�^��[�#Q[u���N�d����H�Xn��#���gp�d>y��y�� �9��-�d�2d	���W.`��x�0��o�&Nk��xb�L����O�\i�gL �}��K2��� �c�g>��KKh��70M=Tr�1�8�Hq�AX�vr��* З0n�G!��'��<o/���u�*@զ��HXȎ��n���]j�f76�U�p�"�.t���̘� �(�Uz(���D��l%&т�>��8�z�U����Ҷ�S�X_�����$w �dft:�Oi��B��s��E&�xq���2>�dW<��A|���6/s����p{�Aւ��sd�
�0\ܪdDb�:��}É������nd�g'p�.�jɈ����)�}�.��������z<��>O@\bxI
��{bF�&�7u%a�1����7���:4Z:ً	J'�s���Zo���-i�m��Y�T���׫�Me��I΅�`|��ա�\��{ߜ1�r��#�U�����W|.�U�i�� �(J�w~�"ܳZ�E��w5�A�候�n=���[3TF���=Rv�� ����
�9��5� �;p���uڦ��c�Z��U�t�VSL�5��c���R_ }Zd�Z|��������;i���s��@U�r�~g@���/a6�;�cQ��s0G�Àւ�����R%�g��.]��Ĩ�����|8Dc �+��P>�*��F���˖��Gt���!۸f?˖*��ب
F��	��:AV�������_��O��kB@9�C���BE��K/(@XZ���A���mki���8?h�sLH>��Y(6�` ��8�s$�0*�5�rTe7]GY	[�Q��������w���/�7͟6�X*�ǷӳcQ��2H�g��>��v���k{5l�e-G� �B�������W��H������*����m���^�r�G���s�}.Mm�uM�=4�ǫ;��eK��Dqq܇����SLC����
VV�k��i��H7�C�7��o5�V��P?в�Ngx��1]lL�ph��>"Qsv��1����v�0����G]��S�����Q�K���ʴf�	���&��z�z�k S
U�Y%�h���S�W�ѤR�o��`��VN��� Vj��t���a�
�l_���B	Ʌ���g��pY)I���t���x�\�j��1R�x��K���7��ggL�6�]�v'��E��+}jʷ.�_�a�J���%�vԉ�S7�ȳ2,��?mþ ��g*��|h��8f>	�ٕ=-��N�)z�,�;��y���Q�4�^9��B	y�b�����#Q�Gף��D>yڅ�8�NR+�Rr�@�D��r!T�����~�Ӯ9��$�V8x�ܛF5�O�.��
�M5��K*���˻���W���`;m�r�HdP���ծ�x�@�e1�9W�8�Ta �L�ֹ#�G���Շ=9�0���ڼ��P\��iѷ�-�>�3��͓:SwzVR.}%���ww��q��Y��4,}M2L��|����uE���Bb���@�4@�]ҁ�m��ma�g	��������C���C���`o$�վ[�Г��ؑ�M�q�Rg�#�'�LU�t��]{ "1���wKW/�;���C���m�aiQ޴Q���Q�.d�>b�ZCc��H5:a�.k�G���zp�54B�֞K�H�*�������=?�Eİ��wE�
`_�K�Wdē�=�ʃ�-�
[H+MYZL�(CFM �T�����e�	�`�Z�R�b�Q�ҡ�ìY&}:M���˟�[�y(kz��u�Lbf�iޠ��Ǝ��
�'�Y�<�	4�d���Ѷ& I�cXJ"D��,kP���iJ!j����/�Z4i����`[|�����U���	����⮑�Hb3�ߪ�>&�ޤa����<Px����m0� ڿ�j%	����ҏ��W��x�b�����s����q��2�Rm@21�5���Q)Q�X�c�sp]%�=!�}��L-���.�pKxM��-L�v6|�C��Zih4G!t
�r��v҉�)�������,@��i��o�����0��r���k7��S5����9��0<�zj���`y+d�g����-�σQ+��G��\�	���^��"��+�8��<���� y��A%�E�k�2_ؕ��?.�=�Ά��3��d������3U�;��P�x8�P�`j��g��}�՘Y캘V@l2����<�9�[-ݱF` N1A����C2��>����58��?�������L �54�#2��C)�0.�X��F�h�vؼ&�z�x�L���;ߩ���VRzi_�62Mv�)��LѴ�u��H0�K�H�S�u�0�>2�$�Ni���A�3Nx5�q(頗s�f$8��ǜ2���t��VB��5�O	����3����r�t[���*�Zi�<�]�L34F� S��o����������/ٕ�=�K�g�|�	y'�7�t���K�+�EF\bל=e�snJθ�b�m��3NR#�I�{H����ڸ��W���s��y�^��J�e��`�d�cS����$�	��	�)\s�(ԟVrxS]�?�w9_y�\�,UZ��Js��g"if��ͣ�f^U.���f�ҥ%���&�0��",���`���9�츟*�u]
�f����2�q�����v�X�0o�F�p�B�#=b8}VX�5�w�M)��z,�E�-3�8q���Fm����(��#�����̂���M�o�Q�%��E�F��c�b�����d�6�R �֔��[U���v�K��S�s96&u!��l;��@�Et�h����O?�\�D��ǭ�?�OdL�w���a�%O�%�6߷��{K��ŀ�\��m7|E�EG�
��8,��-�4!�H�N��b��H�kNa��Q� ��f�\AR�\�0�ɤ�%��2��^�l^²�x��~Z���z�7Չ�l!��)�JQ�}�-���/�	��'7(�ω������6��:l�E"/���|��[~�GH~o�"8"����n	ۛje+?U��]ӌ�Ƒ� }��zz��4�X8�U l&�G?<$�����U{L�X%�u��ň��cI!����`؛��1�x,�"�mo}�5p��@�p��V��V���K�dU�l��G���S��ֽ��E<@�g[GUpe�)i�וyn�DY&Q�a@h�L�Q��}�7�蜉��}E0�b�b�Io�,1�&x�o�?���3��j~�eC[!�]��T�����3s��Ӻׁ�\ٴ��Ⅵ`!#[Y]g���;��Y<z�=.�(�L0e<בg����5���9s}���+�	-��z_��k2d�����Jou����E],��r+w?�"8������HK��� �\6��F�ݠ�"��m�0wF�s��W�^���鉈�S��L�"�[/�A���,� ��jˀ��N�d����aA����ր?vB����I��A4�UP:��w��]v.����v<�)���z���N���'H�!o���tFb�^d�3���.p?��Ă_'0~X����#v/e50t ��K�r��i���,d��n����|R���^����� ��f�aj�����5��S۝�� ]�d%-�2'n8K���-#p:��S�<Q�>���׊�f�O7��/��*�J3�-��T(��Lr[b��33S�g�#���>#(f�)Ҹ+UX�*F��Lzd|`L�)}J�� �c�+nt�_06{�%.j�
��t�� x��
��6�Gi��k+6>$��m�4Ŭ�pu�x�,;��q��ߢ�q�P>�,��F�f�|�-�^דg�l�6����h�j�=hk��&�ޗ��f?����+S�͍���wR�"6�r�F���+2P�w!H����Q�$�+�Z�.��SG�M�։H�.�F���`[�%Kn�8Ѯ���M'��A`�C�裍~��II��QYv�YG�!��$�ߖo�n�M?�m���R���o���݀��?�-��@�[�6�����M�՜��=�v6H<�b#m�(��k��V�ϊQ_t^+��ؿ�OE�xȥ햼�|R��^]�uŸ�A6p�x6����o�/V96|�
T/��c�O�tk�����	�L,^�Q�rA7Tf.�1����"���5��\d�ϙU���X�����[q �P.��Zp/;A�h��zc (���+j���H�b���3�0��DZ^�rg,��}� �� �4:�	Q�c?�V�����3���l^�������!¸	����5����̎��.O<���'�%�����������R8hw�����d{Ͱ �EV�l��i�K�$@	.3�:M�)8���4q�^�]�d�� �]�������Pp>����|-�@��(d���:	�7���>}+,��U��۵{f'�qT����V��W����;�U��}�nʄ�e/�=h�n�*�x���Ŏ�'��rM9^٩�$~'M���ј8� s(��`.ի����W�,�埈�L���U��w���/j���S?�#�q��)c:M������D��WZ�-0l��R�~5���y���v4�.5�/򷝜�(`w�X��;�8'�|�Q1����v`�2d��-�?�pi�����a5b��[��Y��t1�c}+�Pu5��A�Y%c�t2�Q���'�ʞ���w"=����bd#΁��3�f�]-���R��9�/-�;�����	0N_��� Di�c�T5Bfo)�.�#Ⱦ��o+�9��v�d��~,����S�<JXGPh�-�M�
�*4+��x$�7A^v�.݅= ��#M����!g�J٘V�yǆ\�n�����W�gɧJ�u%A�X���ZiQ����cJr^���͡��|-x�Nm�����,�����+6�3�h�F�|*��`� ��#i��#���A�6˾��(�	����Ք��3x�3����V���|$c9�8G �*�&����C�A��Ў߼_Mի72!�b@����d|�o�DE�Gُ1�[�w:��s�9�� �:�����d��t%�J��6M�(̸*-ߗ���'Rǣ�V�Q �e�TBS���{gqZa\�I�.��[d�.���E�I�a�:QGv���z�>T5$��/�w&���<��|xR�a<u.CV���d�*�h�b�53	�F�����? U+�M���$e\�C�I���k���� YGQ|��r��gKv]8G�谮��<}�9\�5Y.��xБҰ:]Y!���~s� i"���\�$�!��G��A��Td�̀tF�?�/��>0K=�#��?0�CR%aN�`�񃧗�M%�էՍ���r�=wQ�j2����h^
~7q������RN��3��A��ʕk�U�{1��TpӛQ$[��Kٳb�YO�/��r�u������S 9��=Io�M?X��r5�O�'��y��=����U�1u���3���H�������8K��b�װ���f��2m)����
A��U�B+����k�!]h��<m�����jg4����͠�;�z}Z�(t�M�� ����z@��jMsV�o�o�N�����:ZN���E�e�Z#<���ff����m�74��u��g
�x�r�h$�Daf����yDg�[QbP(�����/��@hWQ���i証���R�XE#M�`㾐*�j!g��"w�ȕ�����"��q�S��ۖ��Y4*�j�����>�����h㳹�k�m�;�B<��aS��2��m�EL>P��U�
�	���E���<E�u�����gX�\�'X��T�U7��a/˅0���؀���Cr�I�9Ph����T�l���ݤ@=۞�F�o��:;O�X����Ǧ�`	A�͞I;�ӗ ��z��Z�&�?1������r����Tcs.��[�����%v����f�li87��V� �7��H2��9�}�T���/li,R�/�1e2�z�=��h��h<'�E���������b�2ɛ
�jK5e��֍�U���'�1%�E�>�;���� tj�;# ��5'��-�q�����$���}_-ؘ�EDL�}�d �2x?EDL�#z����{@�!ğ��
c�:(�4��~�Q\~�m��F$�i�x�#j4t���[Ԛr`T��o����:RB�6���Q{��=��#|��a�������5���6A�k�8��09Q��s,R��j���bՋ��C���V�|:0x�j־f/�۾��U{Z#��Km�hX
�Ȼ�����bA���ԧ�8q=OX��%g��9%��|�}��'Ğ���Jz�GD3��4�5+�9ž�Ro|��l�-�[K^�-��P�kո����3���G���������ȓ��Ӟܓ7�q�>)h���P�1�#\O�X)W�+.xUs1������LF�;xl�-�	q�ST�_���]��ZЌB���.���Ð�5�Q�?��ֻ�.�@����ܤ�)[�����}E�|j�$�YV,��^ �Cz��F�dk�M��5��8�w�'�l��f�h;���72���\�X��gdZ��I]�	�.2�Q��
7]����	��F�8T��ڮmb+a�?5 :��nx?<�Xx��7���,�^�4IW�d��y�e�Ɠ}3-�����u#���i\�eG���Ӏ��;5�:�:�� ���W`)�_���320gٕ�k=��qZr?�H�;w�S[=% 5���B%��~�=��}�'�aic�$*�&}q�o�	�P姪�0~�)��:p�b��J����g'�r�9�p���������od���7�K���|�y;��wup.����N��Z=���G���w����*���^eXy��3¸��M�?��J�"��Z쿒ȕXQO��
u�G}t [8���=�z����N�����O��'�����l�6dH�p�X�eᛯ;�ύ��~���:?��T5m{wb�8YPgS�V�秈������Z�r2#.r�A
����L@���s��3π�s�_2F�Sx�w��=�"�ڧ� ����5{$��T�&�(�L.�Rb㊞ב��Yq՟Ｐ̭�R$y,���5�J["�ZdsQH�q4w�W?*^r�F�⣜	n�e�\F,|b���j��n|��m3o��e3�:�B~�Ճ�o��E��1|�bA	����G�����;h��0D&2����`ly�a����%��u۩�����dTŸ�^�������.�O�N�2_�x%�#�+7a!�i��;�g��I����2aV���]����v9Fp�6����P���-ts�-?H�;Y����x�������"�\]��&Lʐz�:pI����3A�L�6&��DW��o�s���5��{�yS��º���8��@R!�ǫۢ]k�[��ע�C��z$J�o�Y'K�|=ț�rk57�!=�gi�"g)E���9��Q`Fҗ�"�[}%w�����q�Qm���� ��[O/}�́<@F)���s7D�S]N�^�R*��c���
Պ�OO�D���e���t��>�� �s�����W��5�ŦFF ϲ�$'�V�b�9F.J
�Z*�g;��{Q7Y�̡ͦ,i���#sTs�5���c��[����x��ս?��~v2�i��]|�����q+3@�4�$O\X)Ȫ��nb���{��SΘ3���O���j�dAȀ�S91 ���!����ԡ�b'S32oc׵ibA��g����i�I���
���F�h᝜L4NzM`�C�2"��J�HF~�"d��ͨ��>��D8Woj���+766��~���A~hU~n�]XEd�<gJn[���5y�������#��_2V�,}M��Z�����B��X3uC���\f��xӈ!�B�{aO��w��D�sW���6�E3�zyRC*)LXT=��0}����_+�<Ad.����B�5,��B�D�P@���si�~>hjIN�YNK�TG�K,(��%؍��vN��jtr�/����j��ZdR]7����Ҍ�I1���:ܣ�p�l����M��j��p�P�[:��r����_2z�?T��wi��uh�/jj5?���w�23���X"«_L��� )�J��m�v����ˀ�D�
�a�{�����ڙ����NQ]N+=���#I@�۱��Da�ܙ�L�`sW���rg������K�����~��� ����e^�P���zA������^q��vQ��ʐb�
��{��(Xd��9�M<����������б�'�Fh���G�K���NH��x�YcU�h��Y��:96���X�~�!�Bltm�� k�v�"�?���*�ݱ�ފ7��c)�����U�f&#�	�+�<o������otYQ[��;92�3��Ogjύ/]6,d�4��~4�TfA��N�)$�o?O�ƭ��!R�6w<G�k�\V��z�p�ƈ��)��E��>[	z��W+����KhU�9n��<��R��o�43��-��u��3��jc@S�H��@��\���qU��;��\~�n3����wA �q=I�2�lC�R�J���,��!��%�m�TF��T��!�#2���bݢ��WwP�q��ew��k��z������Q��ர�����\qv;�+ Ҏ�O���6,�zo�w���h�N��ȱ�<��O�6K<ƝW+�̯j���� �M��&�	v	�DX�s�tr�Œ����]�����껮�?S�SpM��{>c�TB�h�_ϛ����C'bQT�`�*	�i®C�ۻ�A kP:r:b���$E3�v�ܝ��=��H�z�C+�]j�^�0d�I0$�f?0:\�������{�v*;\��g��� 6�`��J�+�6��v��ǔ�X\/0v֍ �S��O�2�r8OZ��	����z�p��]�w����*P�Qdz�둷�T�X[�z:}�*�2�E�o���H	=X��ձD� �u�W�n����n��sZ��?1O2�j��8���>d3�Լ�c�}�U�S	��KQN��rC��ȠMp	�,�c��΍��b�>������k���}f��).^/�~a�_%��������3^E1B�ob����۞�E���3a����Hk3�z`�ĉ�@��0��6�3�\1����r��7��$���Y�'��6�u�+fi��@�,��&�o���F}&���� ���0/_��O�]��4f�ឮ����SIQh�z(h
V��kqKU�
���c8�혫�~��"��������9T�)��!!"#=j�^�>I���n�!��#�����$��b��|�H�Y.�e��|w�ma~Z������s*!=w�9�m�S������.��ƾu|f��A��<�c�*79��_����x��B�LS�O�o�ֶ��"z|�����s��I��*I�絛���/�L�Wޚ��-�#@�ƾ���!��˳g��wiBW2�t�ms��|T���c]�T;6N�\��L����Q�N3����z�@Ġ�����a���Y3�JI�^?��$�V�9ǲ >�>���O�N�X;�z��4,d-C"M�8�l��޷D��6&�� ���o�ȫ"�(�Dx�|��')6���������8�;�\QC��2$��ı�Kڍ����L�fF��A����&��06E�5UYm����h��J��c���'fM��A��xK^3&	~�����Y�D�['�6��TN�%NB�)�y����r��5����
���b��.�,j6uJ%HX�tU7I��I>�£r�24�D�sf@�Ş5�R9T���$��<Ag�h� .}�y���M�b�J�v�6,wE�P���ܯ☄�핒�׉����P=䆍�L�c�޸_]�Hiǁ�K�W�U���XN)��Ms�,c>4!~N��Ԣ;�:�{�Z��򬂩>ਗ਼~�֣�*�s��U�6[D�?�ܳ�t�+�f�@|�s�����<�" ��%�����S�MFw��Lrx�]+V&��@�(Q��P}��'!�#ߜ or��ۤ�w�W�w��d�:qH�!���;`P��^c�u���'?u|u��ITD���ܡ��CQѓ]}~����`f�#���� �|������S�����C%�n+��$�F>95����.�2�c�� �@^���	/8k�N�W�we]{^[ߒb<fσ�X�>1���&��l��@���,�U aFW/0͡F�x�� �>��y*g��co�M��$�va��#s�$��UB`�Us㒌��x�Y�(����E�3�QP��԰	b���xHA7~R�q���N%}|�f�N��I������KJR�9�2�W��
-1�{�݋�Vh����<7�O�����^C$%t����J��o�G���VM���d��fUNø��*4�l�����RvZ��^��_�/������h~�Rod��怉�uנ
����<�bW6���Z�}��d�#I�?�Mf
q��6҅�XZ�|x���Y����z$&I��Qn��]>x�ǆ��y��ݷ��&��\#�#߮v
8�c=��G�?Ut����T(�i��XB�!0��Z�3���r
��oc@&4)��tR��;i�k�S>c����歳�y���1T*����BN{gzU#'��R�Ę|P-U}��h�	ևC�u�B��Qc�e`Y��܉������<c�I����H���$7J���y�����t��4���E3��۸�!���Y�UZ��C(%�Aƣ<��mp޴Y�yU��v��j�_s9���q:?�L��\Z��g��B53Y�Sl������
_0�;ib����M���&�ް o�z����MX��1F�q��|����윏��
2�A���׵�*�Թ��&(K$қ�ș�F�ٙ��{t5�_�X�T*O����4��#��?���������=�S���a����7��_���0���&Y�*7�V���i��7-��6�����-��n��F缟�Y��?�c�C���$�\�z��0J�%���%���`qpT��V�>�d�DY�Ͳ�ǭ_sA�Ϳk�t��F%�l���S�=a.�1\4�T����O��)����s�H⏢`���:Ʌ��{w�ϔs[�BB%l��ׁW�`Җ��jb�/oѶ�oe$�M�ċ�!(m�$����L����7[�c=X�4Â��=k�!
Ο�#a*~�;�t,_��(����,�p�t����D~f��p�V�ֺg�2y8�K����k��s�9��zY%�=�f����?kD�*��Z�Г����p>��]�wn��z"x�N��f�T�\��f����G���SALt߽d�L��V�.<�'񂡰@�]ͿTO�FN��)��l���f���E-��|�AC�0R�k��$������g��p#�������l7�O?��������]|��%�-�(/_�LKt�̒mE�T�@y��g�锲捩��ӛwh��@X�V�F�i�"��m�Tt��"u�6,���x�HR8w��W��^�`���⠮`Daٱ�͋���#���Ū,w�3j���w�.��A���JJ�dp;�zG�ɉ`��|�a��3ҷ�C
� N�����u�m�Q�q2p�_�3?� y	�G�6���^��eN��rIWM]СIuz���#;�f�-�>ja#q11��<�t�������riJ�V��1�C��<mp!��!.���E'g�:��YY�$W��&r�4ԏ�f�4঵(�?U(�8`���IaK�R�=��Ʃ��ja�*�#�e�>�Uڍ���$�Ţlv����E�9�Y�.O�D�л�p��Cs�ݚ<�Q�+��H�$���zUEl�AK��푞�ʍ�V�"�������g�t9�v�%�r{5á��w�i1�q�z���.Hצ5t�h"*/t3{��_%TOֽq9���$���n�k�T,�u�[(��&�4_
�`GO�`)�1�l�vMY�/5Oa{�ߎv���V|Zڢԛ���V�cr���������':��oJg�X{F�Ώ�9���~��r��|�@�0�";��#~`wa�ܓI�kPA~R��S�����9�>�7�/�\\�x4�t��*H_M��b*~b�u�yJJ�$���ˌ��N�q5 �9��(�'��o�#�@�;hbr�{��X�q��'�4���s+ST7@~��1�ɫ��`a=�A8sĠ������F��J��Wa_��{w��T�i�H*�!q���]с���q�P6�r����wO�V.�]c?�֭LX�2Tm�t�ŉ�~�����8��B���g���Q�WTV�`��t�ri��N`i���2ir|T{eT�B�k�����J��UC��/������}��5f�V��I��>�T�,��
4Z���Y�&��7]&�
��"f�������&��t*��	U{���������0�w��bavJ0���d�B���I�{;��T�p�9�^�9�D ����T����w�Mh'ܰS��0�);(�l��ha��<�@.����S`[c���w��{>b��f��a�3E���+�;�RHKbN�`�:���/���M��^R�#�J�k���we�`��',�������	"qL\�16�#�����Ӳ��UQ}��B����� ����]� Z��e���qc�)=����U
mRU2�w@C�_i'��;F� �a����,V�,�X�J�S����l��K���of��Ji7\m�"�#u��o��W��uG>"K2)3�/�t�v���[D��;�>TK���!�Hp}�&���������N9= �m"Wq��b� I�w{�y!�F�ب��s��w{JS�ǆ�!�Lfu��Q��n귅,�@��at�-�y�`|��!
�e^�S���&�o�%MM����~�r3dV��r=�)eb�3F���}\��D���Y�yQ�@滯��Lo���H�����Fx���.gZ͆����W�4����ޠ���<Xfc��E�9���JƆ��.�E� ���ޜ��Ɋ�t�e�ڪ}+���\a�7懶D�Y@G{��vej`�9t��m
qd�v�9��Ò�T��N�2�����R���x��nj3�@p�>	V�Z���&k�����N���|�L~]Xߗ:a9��#������gT>�P�C�M�#:չ�I�#��>�P{�9�g#���r%�+u��+Uu=`�����*��Q��P/T�Ղ�O��M^.$n�:��� �X��{��aW+�r�� �����o0cPߙ��KeW���̡=��%F���^�_3��,'�M	m!4���u������t-�h�=;��[^�&���71��y�_e�B?�)'�o2�Y5wz��2