��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_��Zjwެ3�PT��uכ�}
~��DR���I��А�e����+�t�d[����!��p�� �n(U��
W=�O��,��0�L��[p�U��h'U$� �g(��>α�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P��8�t6ll�
/�v�4ei�VD�i@7l�����Y���'_L2�"���1��%�;t��%��է���j�wr�(t�vEW���؍���|����t��	��G �3N�K�L6��K�Uƪn��|2�i�ŪC�d�'��y�G��V%44�>�z�][姴�S���&ZwT��ÃR���!�w�S<����rW��"/�g�f~�i���)!*���7��K��H����R�JU��x���R�}��,�}e��E1��u�@:�zPItn%P%@�Ok_��z��`���-RȎ�z�<p�T���w-c-5��ΉX�⢗��wcI���^c��N~}My�S��[{m\�:�Uɶ�,�Y��a}�=����%�r��
m7�H˲>���U���v�}���}	�L6������8�*�# �3_=0��cQ���O]V�S����az2W�:�/@|�g�o���t#HO�%�=�$���3�I�XlK�[��'�%aH����>q5�\��Oҍ�CYHQ��dT�$�'����l�D�-ʹ��E�7`��g���.��\g�]�̀*��M��QO{�7hN�&���7�6?Y�}��߆��� �{2���1-혖$���r���a�;��b,���ܬT0L����7��E%��	9��}meHWPؖL�1�����e2O~Z���M^��@k�|�|&f^sv��s��n���`�G�CS���o�i.վ�������B�$Jc �,c��a�9�S:�=e�F�~���ȐVn������� /�n@��Pr�5���t�dc���/�M�,�����dG�[ ����/P�٠Ue��͉�0�7�;����c%�U�bF�ѷ�cOg�_�o1��=
E*/&�3���
�Aa>�k{Ô���,j��k/�Ҕb�?�nf����
~i�G��ԃ�gW�ABnԱ�8����V��J[.�w̰���v��cZ�B�(����π4t�G��S'�vwz�U^�ӏ�1��罸m5S�pM������S� r��Zv�[�gfp�����a+�d�����8����z'J&f�9��9�p�6�A�T!���oמ:����1
V�pbCΘ_Cp%,Fޏ��x��(^)��L�K�9Y��jc�sw�����%����u�w�u�˅Q
���(�og�p�P�%�6'w�M5Wy,,)�'�G�iE�'�I����V�s��ч�~M2��g��ƌ�?˙�w4y��*mf�P���ЎBG�K�|s�Y��ح�{�Z.��Z�P>�S.��U�=�3eE`�-��(,�߁�?�,3vyj�T��Lҿ#�|��u�ո�X{w�h��*�.��- !�x|Ƙ6�f�g�=�n��X'°�ph͓��"���W��k��*G�H�M��U@(�s7����t6����=rH�I��zy�>ǘ"Y���+�l��I�(����+:���Q��M4�!9�&|)���$��-`RO��=�1⽫MO����M�cB��Ј���h�˱Q�.^ձ�_��CUV2�g�0����L[��k�.x�XW�=�V��Q�wŉE��Y��{���S�M]'��׎�)�o�Yki;i�\�b���G_����V�����X���.�����S�0�1=������ l���,-�HYZFH�����3@�]�kA�ľ�>[�9hڣ�"���U74��z��C^�~�J�cuEj�F-@��+|o�ybX<?�x�j����a~q#����M�;�z8�]JN����� u���&�S��N��1LF�	.�L��o�i���s��ͅaF���o��W;:�3�B��=Ju7V!WW4DP����V���Xji�����[�,�6f|���/fL]X��tT�h�}�leB����=�Y<]}`�T��7�& ����?�6~�0�����a!���P7������t��&QClmڱm��n�Gt/������AO�@>w�A�1�	�-�Hy��;�)����I�
P��U2򰆥σ��������X���\)5��km�`�G&J�Տ��?JPV@L�~25�����yԕI �F�/�y�-?e$Ծm�G��;��B� ��&�"=���P�����rC�R ��ψg�H>�_�:�`I��� �A^�R�bP��d�*(eJ��P.���ɲ�D�B����O��b�)�$�?μ;�q{A�������&y��f�3���j��i�(�5@<��pN%=��� �x�7�	0����^+R���|R��N�����T���I9��Fz��{e��0�͈@vnh�2L��=�.�Y�{W��B?n�\�7�E��i<�>���'ڤ��^���C ]'@e&��w�=�:�-��&��zpMyɄF4@;&���������_�g��ȡi;Un�%��\�q�������k�M�Y�Z8X��`{�5��s1=]W�z��˼��qD\�a9V�t^Ceݵ�;�o��_]�׍��y�2���X��6�x^��	v�=�����`щl��N&��n��nm��yL������o� X��C�XW�3��:�=��ʆxj�����_-o��4 �a�����>Z��3�-�
�+z�{O�kbW���ɸ����z�Q&�t�i>+�ڄe�ѣ�T���蜯/�����BF�q��1hpdh���
�q�wb��^_�����Zg�л
׼����o`�
�%SUOӠ��S����3�����4[����;/��hiHC�܈��練�-dj<�o�+�o�Oʬ��5`6Դ5��q��u�E�$#�z�fm��������!9����O��驳}bw��:n��QZ��;�DT�m}\�^>���AZy�/�XZS9����9����ϒ�\��z�:��
.$l]������"���J&�>i��u����͉g'y�=%���j]_�k��j�Ah� �ސ��␑n�Kv��Fp)���"_���ȓ������f���v��J�zR���fˆ������l�N��u$�IE��#���n�+I�n[bI���y��B.C�=]�0%	0�c�4ɚ۬Mɰ�ӕ�~A���ӣ�ǎ��Y���$�L���&��h�VԼ��29��aZ�}ڒ�Ĩ������Eh�T�o���yY�ٻ��O��V��<�v���h^(��	ll��;��p���o:��"��BJI����I�}�	�'��t$ʀ�]���jk��́�e�{Q��q��R�F��gD�W�=��R}�Q7����^0��f����=�$�m������a+�:���Hd�&�H���M��iƤw:bs��5��fSp���.l2k���j u�$���� IqD+���QΞ��w���`�\��:EV��;N_�s8D\�V]� Y�ǥ�^�}�����}犴�5���� �e�D����)ԧ\簴�
{u�̹��Bo�(X$��2S�2��5��V�����Ʃ/�1G~�3M��e".^���]���d���`>��E��f���'r^�;p$�B��0a&b.�Qw#bl��N��RV����h �m���o���ծ^:�{n�r~�N�u�*���9#񸐗���O�8� `r �m�>n���8��_dt��M�7GH���t�
t���ymMh�Iv���/y��OE�C�6�Z�E����|��a��|H/����O5���H	���}uجckXR1M�1��
ِѹA��̒�n�zS� ���&��Uϻ��׽�)1r�ʢvӗ����"��`�ޞ�Ã��=�)~-���#�Z���_�Q�B�Y�Xy�/OBea�Z�~�dқ[���$ע�'�/��a�L��#+�[�|���7�t���P~$�X�{��&.���J��mp	�h��~�A,jDo6%� �N���|t~�]�=��Z��ͭQ�$:A60&k�ׅ7%�7�N��7ѫjP���Zc�Ŀ9�9�*O�1�����u`�#$ڣZOlwџ����k�5�rׇ�颅s�7,\��a�Rp�f��;�l8�-�����3��K������!ZD�v5�O���VL�'�Y�pT�����-0�'5�U���2ᤲx�� �,H����Cͬ��9��+��'��Ud���y3aP6� K.�ǯdp�'�m���_�(k�o���A),�����U7ࣳ���@�v��i��_���>�&l�W� �F��� ���F�:��7�3*��
�<@-��8ǗX�K��҅�5�&�����*J{d�a�:ϊ��~@e`�:�]��@���J�I���DJ�e�5�Hj��=j .�j�ѷ/��j ��]gU$O:]����|����!:�R,������0�$I���=ݬt7�x|�����>AM�N���?���蔈�$���)|[D�ps}X�D��'-��I�[ue�½�P��Mp�{���&h]�&�˒��m��al�L��)�s��vpW2�X�V�ygE�\(~��2<�LPA��	O������X��:M���o�:Db͟=���G ����)��h(���o@����yhh�%H���A)��5� 3T��m1Np��Ha��H];�;��������"+*�U�^Yv�Ud�O���\�s���J��fT���o'���\��+���l~�bB-^�
�J��|�a�Xț���c t��
�OzWw�]wjB�빼,$ܴ(;n�Dau����o�L�$�߶��S��+j�<����!h'j�+悶��^�Ɩ(�;&�����7�N?�{��VB��4����lFp�z�E�0��}x�o)�g�W�_����z;iº��b�X�-��uF�f=q��? N8��H:hC�������n��VGvY� ���h�f�n؆��`{؉%G��b���r}�R�Y�t��W��^��.���h%���h-Rϋ���O��5�!�.��伉��ޡ�q�+�lF��^��dQ�$�>��F�;���v��Fq���ÆN���M:�J�D��ˌI$�e�Y ���Բda����R�P�|�m�b��"�sY�R�9������@��叝��~�Cxf��&�Pd�������-a�U��챖
�m�t���a�x��m>*/�Dfy*Gj��l�-wM_�Ox]0>�R��e��?��E����[��\��v�L�Q��8�i�Ŏs��ֿvCc�j!��o��1H҈��BQI��@�,��¯��rD�Q1t�eM� �V�����f�-���x4+'GEy�-��ASn�y�����Nt���l@�z��^ā��q�pɥj	�I�hJ Q���^�����R ~��d�O� Fm��;�*��ג9&�2�&�4�m��<k[�j&=�����p"��R�P��Iz�QzSX��[P��QT�Ւ�;����<Y��/�2�p�<)By�(99�/Ф�����K0Ѓ����|��>�zg3� ��dDi._/��������>K�Ez�0��uf��� ����\R�[��Nԓ�Z%�'Q��cGtg�K��;�#TW��-��R��kg���Ef[�HFԇE���f�q�,�^"���n�C ڊ.��}�9<�b��m�>�����.�ln��V�M��rH�>��Vj�/6�?+��ƒ�������f����DBϬ������6NǊ%U��qU}��T®��x5�7$��Y#E���+�ɩ�=��ـ0U���d|��C1�m���@0�F;�gE=�V����W�nԂ�FYz��W�\/�2��lJ�{R��V�����:�ȓ����ȯ\�S�7v�w=��c*"�l��H��+������L�N�zng}wZ��o��q���n��uM�a�P�w#��K�����:hkh �m��T�y��5���.T�Ԁ&�d�g�1�d��w��0zR���]+R� B����Ŏ�	�\�~�p\;DZ��>�K��e���^�C6�����K����QΩ�n���!�\|[W��v�I2AL@�LٹKp��WkA�߫�
_����B��Oi�!��Q���ќ�V=i�#�O� 9!bV݇�X~7D��AS�S����ɜQ�D����1@+{}�:�NX��ϟkB���Lu��8�c��X@OJ����K@���`*C��t� �-�e�@O�w�t�i�n�K��ι���l1(���x|9g|$��iw6^n=_o��[`j��]t���01�_#��EEZo�r�<�dƹ��;��l�  �!˕p9�H��� 4�q���&ӿ����N��I%`�N��a�vzJE[fF:�c8&#��o����z��:e0�)�ȺƆ�e��C^9w��:�3�|�_��0��#E���~��������[�ڑ;�Ȃ��Q��0���-t�1c�s�6:�쉑����ř	GFP��!{��w��a�	wd����H��O]��?�S�!��&c!�|k�.�RV&!���dm�E�2Eg�M̺�����`c �:E.����bBՄ��s�ɨP?����s�D3�|��ďT� �Ty����4(���0/Ti�M��uI	zO�Q��M��j��/��a�[/����z����h���A�s�+�K����u��H�EӢ5�8�F$ʕ���m����h��ԟa(�e���~MU|"	�x(��J�o�Oc}u�BH媹��`� �N8s=b=�q���V#d���V��;4^�C�@�X>6i���?���ai�-ҭ�D�eL�wT��	��u�K�Oo��V���b���!�� �i^��K��h��PX�yRH��x��@.�;3�q���MV�H�z�*�]0���JR�Lh�o\�����>J;O�چJ�ɶڨ���ŧ=�^)��.��i�V� ?4H\>�l)z(w\�T���/Ĩ̛�<G����^���@���O?d�-��o��L�Q_����;)z�IĲ�^�X\�����6�%���)����gh!?�L�!�E�,��EC�3��W*�z������U(�����.��]:#҅D^O��C�J᭥���e �x�t�89R�[��/�Ea��m�/~8fF�L�cW�~��ڗ�?���T_�1vv�ٖ���C� �#S�����?���qs$���L�"��e�ڔd��xj�\h�(��o�"R��Jq���tK6:�+%vc��A�\����ڗ;�H���~�EmVДV������u�J���'��3�Y��!�X�g�m�Z��EFf��,����_x1Ǜ9ηiy47��mG���d�ͫnB�g:��N��7S.�o���wx�Rj7:.�4�!�|�)N�^.�S��"v5��f��6�����9:3��ɾ����;��+�	r(�������9�Y���==�ȑ��Q�O�������Y�h��^r*���8L%͜�M˟c���N˛+.��L�Y	I�>��'tf!-��3��6�K��%L3	O���k��Qz�V� ���V�,Q�͑{E3Hh$|h����AX3*���V��3Z�3as����
5-��C�%�:��0p`Z�=�2�yh3�C�M�!�v_�m&v��l�\��|�)y�I�a�o��N�D�������OĠ`��II�E��_Q��R���->�j.�f���У�Z�5��u�F�>�	=������.G��n}"qC�w��:o��/Mi�L����K)�����u���+J��m���zqtw�b������8=���C�>��S���X�F�PS �r<����+�O͕Li)�@�U���9�(�����ҞJT�>��[� >!�_��$�ft�2/Qk����Z.Gb�� (��=}_C�]���J'�v�/��JF���-k_���
��#����Sс�e"W�!oľH�x���W?{����5e��N{��qQ� ��rG��s�Z�ߙ����ũ����dl�QS;鮌�	�������6t\�q*��b�o�T��<df�+#��鮃l���j����N'+D�z�eW��}X����š���&���sC�D��[:��
�Q
Z���33�%�'=��{��V�o0�N_�tZ
�ޑ��f��a���WU���%�9hq�ڎ���Gd9R�/GT�s��Vgy��Zj��<j��!�j�w�_���;X��ğA�b������ZNO��a���>��@d@�Y��P�R�F�$@�ܵMcqY&k��2 ܓ�ޫ�=i�9�����D����ƈ���?7�eᨑz��4(��
����;<�g@v�����&��=V�����]�b�H���tY���ҷ�ԓ1O��F)*Q����S[a�;�X����+{����QI�T7��wO�_�㌂m�`%zU�ֳgC�C.�u�֟M���:��y�8�t�x�,2o�j�$�)9ڿ��#)=�#Ļ�KW�,�jH�:V�a�U��`:!qFB[o������j�2ϗ�U�)I�{;b����h��n�jP���i�0�`����p��j[Ѭ����N��?]�$�:�)�p�c5�4`�ɕ�/�s
P±y�S�sg�FY�^�<��q��5U�6C�(lY��W3;�Mb�k��������-�X��+��B�Qg�,�J�lt�w�q�����Lq-W6����4J�����s'_ �xW~���	��[�:\���lN@H \@��p;I톋R5q?�''��ӭ/j��36�����6-JF��J\��3�Y��/�$	�=��@ �5p��V��k��Ռ:_��6��lM6H>�Ӊ���wEk�ؘqf���ǳ'��$��2d�L���,C�3|�қ�k�Y}����-���:�H������u%b�`Q��m�Y�s]׽��6�����c�����,�|�m�n7"S��`\�_�=�����FY�W��sQ04�Umu���X���Q�jLc����{4bTb�ۖQ��ѱ���Riab�Yx@�4�!�#x�67�Cs`b�#����|c�d4R���x�'��L_ ��D?�PE9����'D�{rҰ������`oN��}l>��� (�v�������&�O�fN��Q�q!_:�©�'�~�4NR�(�h�dH�[���s��ܫ��C mC�ă �[�B��T���r$�n�UpP��iن-K���m�tO�B
j�pW����ߥ�wY��Vz�a��|�������Ŵ�_��ڇy	=���߅�	�ga��f�n�0�Σ"����h���"�����`9ƾ��.�8��j`.�T�~9�y�\D�gZ�%
�؋Ĩ�-V��PRE�t����h��T��w؝�nK>$j�>v�Z����Q�|�0)k�}brf��YN0
��L���MMsʸڢ���5k�ȓu�d��/yY��]�ē��8��Vx͑he(۪�t������������M��->ǲO�������#��_BX�c�ε6 B��`�;����*��&)�����0oaN�E��Xl���%6�9/�Ho�5����ș�7iIT��Z(��˛r��^�'�,9}G��[��3m���H��ƚ�`��I+G�����^�)� 1A�tY�@��V�i�qRH@�T���T]Q���d�mM��NP���ӓ����i��=Rі	������DC��������%N����&��������J��(�g8l���'��D�H	��(pk,����\q=F�<`��� ���ꇐ�!���E�ψc��]�]g�	P>|�P*��0>=���J�E�_�TH=_Vo >B�ga�>�{f���elK���j���Njʁ��}Kd�g`I�-�)BS�h]E���լ�4�aJW�iW7�~t�0��#W{Ǒ�j�Y@��+�7o'"��'�
kli�L��e�����R��_2���8W�׺��k_~�r�����	���I��~4Qb��q	�F/o����
G�)�n\�N`#4�(���< ���������R��&��MU\gJ志���j��"�� Y�{�)�*�_���N��@�*�.�3U$�T�zy�X���z����	�}����(�h��O�%�C�L�4�Zп����Oy�;C�Q�^�������J��>Dn����X�:��k(�I~<_�>G�rK8,ʋ�]�_6�\���	f�x�7��lծ5C���d]�iP�*��s�"�3�ݲw��{���-tP����W����7��4&c��V�FU����@�j\_�sw[�B�=GO�H���p�q�����4��'^�������/0��55��L�10'q�pq�0��%���O�H�K�F�o״�94��8���hVJ2���̯0�D8��1�0�J���I4�"��7���b���>#�5�i���>�7������P���U��Yh�}@B�f�t��wf�C���j!�1 /�L�_X��y��j��$��ĸ���Ǆ�����2���'v���ƣ��� ��>�5ܘ]�e%Jp�Ԫw{���+���B�E��a�N�����cL��4�V�8�����Ң|�iG)}��/艶/��s��bH6�
���:l����l��$���j��Lrmk��[��tn���ݷ@ P���-ׅ���(���,j��~�@�r�#�o��C�.|�z��-��u�$~%��O�@~�h��E�O����#�s�X�3�ڭ���cB�o�x7'����-B\��2����l�âw�S�1.��'��]��6̌�����E��s+p�j?���y
���s�Z= ��ẹ�H*�J�1�ɫ�a���(�y��]'8�8�~ے���<�L�>�����l��I�{|�hj��ʶb�r�Z��������������4���vݔW��.o���C�oY�D{���<~��3��V�j�/ΙG ����S�ɼC�,��rK`܎��;�n�:5����{�����]rQ�uuN�a,c�����(��uD����ۜ���u^Ͳy���Sх��Ο����|���F!넶XPٟzț�t�5�M;����~��V�N�&��ٹ)�A��JG{��P�f�l'��0F:���a���n+�f���C��|��b8��ڳ�����;o��,�ݓ,\�*ݑ�MH��0h�ZY�, �D*�p�������R��3	�9�Xh���
~ /i���� ��;�hН�Զ�3��s=��H�
�v/XFRA\��w��,�gӻ�V�v'P�R޾�%�N�}M�xMxDGm[,��,|Y�Q)�,p�4�B��#mU�Ӧ��9����ɦ�;;"��ɑGR�Z~�LB�y���T9+O�x�����v1jc����@�6J��D2�y���*�-U(X��]���ҥ�# ��9���wF���c����x��)X�����-x[�ͅ��tlulî����/X�r���(u8��)�����*=��X��j1k(Bc�3H���d���q�Qݍ�;Z�`K$@*+Y�B���8|��ӶC�C���� �o��'���,��{�5?+����)G	ۚ{���g� }ݏ�*_�h{�вB���_��I����4�WT�9��8gK�69jYTxHEG��`!�?(쏟-���zW���Ï�`�
Mq�:3#J,+rل\�2E���10q eK��I�6!��S_��C��lfG�����)7\���'�;\ņSub�.�'�hv�UO�0��6e'���u`۝�|:䚮���%�+���9m{^�BU�[��g����3�bJ�m$,�ᤍye�g���y-"���nȷNqz�ಓ*��R�DvpQ&whӐ�*y�mi�ߏ33@�%u���~��F����t�u9�钐g]4��er?���d@! TN���<Y�ΩZ+����R��օ[_,�iq+F�u�;�3fe�	��=P���Z��c��2<Q���=m��-en�!8��fۍ�9���,ͮg{�9%-� ��'Ҷ�*ŕ,�מ,<��]�6���i4���9(w�d3������b�m)y樽��c��*a6��C�k��n}�����H����8U�Y�ds���V7�� s��݋9]�u��4���^���A���yI�3UvO�M��B�&U!�IL���,2�D��(֮����KS�@�-0�5�')'�'�j�<>6�;��N�ARlIU)�U�p����dS�ӂkte��i�=�]�Q�=rit������R
��}$D�cʉ�=Ba�YCѫ������DZ-�����Ϭm�G�����q���
�|�x�P�w�{I���6�%gԌ-��P{���[>�J}Q�	�N���=3u�(B������GI���L�<z
N5Z�Շy���z�2�^��:�`���z
�ǥv���ϖM��oSZ��O�L���<��u����e LF�^�x��Q��A�}�P	s+pF�Z0��S1ʧ�s�k���N����X@O=1��f�k&�3o�~~���>�8*��>E|UZ�]�Ł*��fO����P�su�].�l��W���į�,}�ݞ�?b��v#��(��Q���;���?�0�t��F�����g��^k��$F$���		��MSX�tD]1Ti�v��-�l�[|ȁ��Rh������C��PV�}��x�����M����p�HA
m�gfP8w�W�eJ�ۂ*�p6^]c�5�N�w�*���Q��`3�P��w�:�j�gAB���'#*0�Q��-&>	5�$]��u��^�Ȱ�F*V��J�{�����z���=��Ke��<����GQ�����NL�{-�/L�I'���g�É�q��f*L��2��cK�^���3��+��"�6oh�k������z髼��>?�5��D���eu}P_�%?�^*Y��?|nT*(P��߬,�(�Ay@�q�������	W���n5'���{��߅�z�r����ta��G��U|0�In/�,O��]~G
��u0dKJ'��v)�5o/��u!��NE���N��|MN0-���$U~*gNF5��jc�0�n^��^�NLj��_�HG2�e�>��Ivcj��_Ĕ[k\��{2��ƾk� �(|��W<�������|MŠT���i�2C,�������'�	K �^�6�YV�JO؂��κ_7Ndj��XF���m��������iX.��b6i'%'��պ����F�h"���5��}2!5��^l����S"��II�g��`�"〻�4�<�Ɲ�an��Po�'?7���� v��'�u�;ڢ:v��� ���]Pwf��902�=������������@���gࣜnJ��y�-�og=��p�JD��f&��r���{DӮ��aSW����*�I0��[�e�\9mAz�&#S\Ɂ��E�Dx�n�4I�H��X��-q�O�s�|��q�n�]��͒/#t���a$�@�1���W�� ��\���Q)��M^Y�y�?9ߥI�h~]O׎Tf���Q�p��n>'�n3V��9/��`�pƗ
uZ�u�o/i;0���*2�:��B��U�,��������2�>�h^�,c{���Q�ô��d!-����[���s���(��`�E@��s�;�u`�4]�>'�� �L�;��(��YRI�{�?Z9�O��д��Q?m���2�MV�D9���i��+KW[B�0�B�j����'��p��!v��(T�#=e�~�&�:��6
��'����X��e}�W
�<%�A�g�[����{_g�G"����۠�ಮ��h����|x�S��d掝`�%s\Í�sF�@�r2����=�a�H%վ>/X��P�H��RgJ@%G3����a�<�K���N5<{�㶃�BN5�z�	 ��P�#�C�V�/:J���E}7�@ϏoM�`�������w�aT�s@|�̀o��`d�Ӽ�]<�|?�U��{����kH�2;4��&3A�=��g���xF����9*K)#�RZq�k6���_��MC��ɤ��'���]�6ٛ%�����~nl�-10K���H� `��|�@%�$!%���L�`��s^$�+n��d΋�Ȝ�.���:p���
2�"0��D`L����b�%�j J�7iB�訤�\gp��'�E��J,��I�[O&:{z����&������6��Rԃ-��M|p�Zv��%���ٰK�� �k���R;�-�n���ؼf�u�֜X׎Q� uaV�r�(�L/*��8 �\�j��� �B4A�Ö#]Շ%��bX��oB���֌�(�.ID.٬�믗�`�.-_�������^\9����G�y����Y�C�i@��[J�|���Ҹ!�k���G�f˸�.����~ҽ�6=���CX	�ԡe���j4�O��d��틤m�w4�x�-�}���ǵ|�0I2P��)�|O1�Fs�PX�`uLc
�/�cy�ɨ$w��I��D�*p� w� �@VUa�g�x�� ̅�φ��٢�5�Agݪ�rR������v�k$�����3v7�'�Y�8h�u��o �0 T;�I+^�H�ذ-�ld���l��	E�I������t�7Q�/&�_,]�qMt�<R�W�K����J����ϑ\��M5�G�J��;i�H��oG��W7>K�+���vS|5�]�,p�˟�B�n�W���Rm��/a�~)���u���qpp�{i|��1��[-�-�<X��Z���_QFϳA�9������,�<o��q�)�!a�	����XI�+)���秢t��FҠ�C2����A˷�Qm}ݖ����R�ӕh���L�n���W���FD�������b\c�T��5�<s��B)-[�H,��c����|W�څ�0�u�um������g��z�Ϊ��(��Q���:�����L�SdF�~,?D/i���w�4�R4�B�9]�tE,{�O}��=ݷJSff�;3�R����a����%@4����95+�fT��!ѓ\Tg;��2�Bm��S2���V�=?�����!�B�|��7Ƒϟ��&�ĭ�W�]�0g�y���EPv@�QUU�:�H@W"�.���uy����5���6�xT!�c��-d�PiB�5�񅋉��Ē?���<��J캅і3X�Hm*�-P��Hջ4�$>a�#&��1�@kx�j� bC�5p$uW���D֐&pĲ�/��O&����,c㒴����#Ǒ
�r���v���|lz�	!��
��yn,|ܢI(-��@Xⳗ��U.�|��+ �wi ���X������D��'Z�f���E�o=���o=����������ۚtm.�+�]d�1��a�	����`*�nZ��i��^����db{�ma�����O�""'��]!>�͗�����J��c~M�GY������/%��"�	����߳
��2�9%��2��`��s���a��,�:̣��e�r,r�����r���Heo�������f1B�9����t��d�g��U��X����X`\	�3�ѱ8^��.
t#�l���I;�����O�n� �;}�*
ᆭ���(�C�ɱ ��v��P�(VH���X�d-�1�2�72fW��9������ٗ�{� �����u��P��ٚ������t��:Q�奇�O��@��jH�y��)*3�M��U,���]�m;M����0�����]�_���|(a�/�6�6�Ʉ�^1� |�u|�	@���r�TK�ݤx�e�-�S�u�R;��־��SN7���mN�DN��LS�̐xy	���тi5�ϱQ*�p�> �2�T�9I�ީd��)h�K�b�v�7��r�͋Sݹj�uw�F��HN�0g�8��I���*���G�ѯpiE3�U����)V��W+�D%m���Fꂐ���Wx��<��&�>�����w�����hF�kq��_/Uj�,����6t[2,,mZ*P�%HZ�o���Zg涯�Z���0茋����R�8#��������c�S
""5����oz�N0��̞�XtVa9� ؽt��jn`Da�3n���Yq�L(����6���xg��\��jN��\eأ��;��'vd�P�4�G�����;�߅�Ɔ�/�y���hY9�e����+ 1/�&^���q+5�2� b�R�t��::��z`S��m8ԩr�9�99_��i#ũ~C���0���*��Ϝ%n���{�� ��\��W�x?�yS�Ա%�-w��@�6�";<dWt���{��e0cWz�� �HWM���U��cc�K����7�3���W�mুG/km��B@�'�!t::pɁf�Az(ͫZ���2׉X����]�I��_�U��"�2?���s��V���	��Ju����#]��|!��;�x�Ň_�=���b�����eig�WV{��i��a	��r��i���I�?cS�/e�h/��x���+�y�,�17P�r6���d?ծ��c>�[��;���?������ڤd������CO��n��Ry�&����;I��ݷ���Z��O[l� �F�����Q�W�X�8�l�~xQ.�W-��Yaqm@c�x-I��k�����
�:wNdrH�S�h���mC�w�j����Ӟ��O�����B�����}�>�*�zvI��L���S�n�kf��*f�M2�n��s�Z6����С��-���$ˠe�3f|aY�U�5���������pKq�$g�b��'�d�ؔ�73y��;mp:��HQi' +=H���#9G�.����p�.�w�(z(�p���u�V2�\h�V�����Hqa��QZ�":-�ŏT��|_��<ɀ�~T��I
mɶ�|��k��2`Y����R]�R�������8���P$_N�-dn_!���\�3��r�lj��@� �F?Mi�1��g>��UR]a�t=���1��!�M5u9����w��#D<t!��q
��l�W攱hF���x�Q��tC�����^J����ؤPjnl�M&��b��
��H?��8��
��#1Ũ]6US��E�?�"T(d�����+Ba`�������-�\�P���FS�h���8��,���`�)��^b�P�'��ǋM�cPN$>�/����}��{Qa V�O�Q{Z��Eiqa�y������2��?�ⴌw5��M�̔
 �0�98_!�䊚 �X�o�P,�
���1M"��8Z8o�y�w{�m-�b(�Z~��I��r���X-���Go㒛�:F�ä�j{�)!�`�����KÖ̒���P��4<��b���U��Y0 g��r6�r���0'E�����[�]m�Gh�6`U�G���\\\\����Va�`5�g1����`p�nc����X��¸��^�$����T�Q%���໵)a�)�������a��@@T��+�\h��q��/ Y�����!G.�R�����]�K����sr��@��+L��}/�{b��ro��������c��� UR�.I��J�
�ڒ��Bq6�Ԅ��3Bt�����K˪^��\�x`��M�Y-s)D1/��4��O��T�iOTHoh����=K. ��.y6��y�Rr6�ۅ �R��1���8q�gJ�vܹ� ��f��Ã��c��� ̷V�O�tP�^]ؙ8�[�$�B�i���I��	����i��Ҏc�������w\D �uw������TQ߀#5Rg�1'�@��.2���k�}fm�&.D�W��u�l�yǾŝV�0|�)���&�(3C>���aE��맧/��v�Ͱ�r��<x�kP�L��\0����#8��Cp<��*X0TG�=O��x?KC/�6�L��e���/����3��,�y�*]u
��}e����n\u�»���6)#�g��ODH���1):̄"cL^�%��q�� _�S	����S���V�I��C��π�<���!T=@�%�|h9�B���0�"��9x�fw��;u���-�OWP@;�8�7�q�x�[��\��;
ӿ���fNӂՌ���AJ�w7��,/[�H5B䰉1����u@����nw%G!8�ԡJE�� )��u�V@uag5�op�PyȶBC�����x��i���&�x�;L�sR`۫w�! �v��QNo��;��F�s�+i0EY��GHkW�f��I�������;}��oν�L�k� Ŧt_ۚ�08�oFrx8
t_�a�����=O�|z���丆ݮ�ӥ�{�5�{�l������)�(E�XUw��<0��������#y�á��?�8��I����{48$C�T�}�rӼr��i�� ߧya]I7�㾴��J3gR��2���=:�v}0�*{�2tf:��}'��K�?�]w�7�0��ӹ͚BBh�bʇ�"���uCt�����~�QBܗ@A�'��7�Z� R�`�9�=k�0QCի�ν'a�	�1���"�����3�7]�ޱ����B|���蹑�%R�7�r���l�̻����^���"��_G:���Z�"�|���\Y�A���f4hΧLֶ�Ts�\�ls���i�S�3��]S�j9H�g�\��+���҂���:7�]'���X��X�9� �ʿk���(T�����}�{�d=ںB���xi�eŔ̔@����RE�~��ImF:�◁��� �i=g��s�p�?��v뗼^��s��AlЌO܂�񩟹��'���s�de���qm�M�������!h�-�PA��>��X1�(>Ӽҡ�n�����^8O[ّC���u�&�,V6���Ee1����ܝ��uŁ	1�~)^���)���~�4��d�#��/��g�UhH��M�\�l�܍j֦�E#⑀��+M�?�Ё�`U���W�D�+7�2\nt��돛��~S�GO׮|������)�_������W����S9n�f�:>$�6$�+�~΁6�g��Q����+"�1^T�P֩��)V��.��y�>��2�1ݲW(��q2����z!d�ZHR������Ge���ү��+��{V��fd� '�$���Ʋ�j�i���k�[�A��YŷSw�b��7�7�Ӻ�ѪH�-��qk1���*�I6v�N�������c���QnI�[��G�N����J�Kɂ)h�p�Kc�W��*�h�px�ω��n�`���sT��R�-e�&�# (�D���u�f�1F<�]�����Hݩ/�&�@�h��r|�U�  � �t{C�7'k��k��%�7��ߡ�]9�|�4��Z1��s�Fm���[ oz�{����	Z�w��״��S4n@��n;����̵�8gM���	�!	WN�[�G^`1s⻻8�aW8�]��,@i���O�v�2�Ε�9&�$��N��-
��T@�:5�j��O��֔�����rȴp����ڷ�(9����4�/ۭ�a>����4f��k��|��ݳR�m9�lD�����P(i�m5�Â�h���`B������chbBphɼ��՘���HV��.Q���uJ���cB��{���/��tϭ!L��a	_��/��'S¶���:ɧ-�$SG�A(�!���h��1��,,TO$oq~��|t�7�jc��kr�2C���)�����t?4tJ<L9���ݘ�c���j����*�)���;`8��X��!�'���'>��dN-[�<ݮ�d)�����L���/�`4�ҩō��H�m��R��>�*p�k���r<��kIC��o}�h8xJ%RJ0˰^���]��{�	k��f�%��f&_��G*pd[C�%��^h��V]?R��	�r?��ل��j��WAu��Z�B���N����n�*_n�����5��Z�W�͎PN�r晆���6|h�n�H�,�k��KqKd3'��g�b5)� �G_��dE��{��)�G���{-Jq4:�8�j�_��/�ήd���=��L�h�:��T�N(�k ͪ��u�}@������.�cd&�Q�W�ǫ�m
')�*��qb�h�}>��!3��u��y�|
�e��� '2Y,��gQ�կ&b1�H����3_�W��j�O�Fy����E)�!�$]�(�aw�@����iʵc�"u�#Q�?�~���N[=��RyfE��X�\3~
b0@&~�1M�<���Q7|VQ��z;�d��������|�M�|.�K�������db����ɩБH+|c�T��?}���U��큓�j�����ڠ%�3U�Y��9�d]*��Q�a����m�BH������e����x�J=ཚ���{UqM�H� @���O1A@����=�c����������I�>%�����u#O�E2�f����z1���gRMC��%q��r�/��0V9u׺���9Zҙ��ۺ�Cty��C� ����}��BUo�1�ُ�ld!/���Ŧ��2�1
"m��p�c9�cI&y�� ��/"m���r�ɪq�ZL�c�)��b��LV���j�@�/F�����6dg%�u�,�K�GZ8ԑ>u��~Y
�B��R<ς��*�4~�B�ss�~r��tlJk꺝lQ5{2�����ha9Jay��e���l������K&�H�-�r�&�J@d�N�j%/~%Ñ?�G�;���9;�a}���Xu���C��4XհU_ʟr�� %Í+�׌��)U2�d7(�������6��Pc�}���\A�0^�!��;L)�x��*��l�2�hV����
<���!|')vFXzK���#u~'7ń��̥�����f�FQO%���1����B��֜�ho8��#/\Q^ag����P����D_�O���Y�$�/�R��YN�щb�2�&��Ļs�:\c�sш.i3���[���^�3���+nj���^�[4��"E>8��B2*~;����qH�	_�Y�B"NG��#�@Pc�Z���ym'��S�S[��/�ͼ]c���g��"���m�b1l�� ��t�@
3����e�U����NG>�Ks�Ic)N���^��|�ȗg,=��􃟟��r���3����`�z���"D��:�'I�K��\��E_���U`��X�`���S��S��=�ɰ�ņr��5��G�=Po
I���(��s�)��Y�ݿ̹m)��>Ҵ'�:÷� �����E�r���+h;Ě�@bU3�Y¹�]N�mj�%ё$Co��dݓ�P�]���`�����ج��U�'a\���<�I)g���g&2����P�m5��W���Ҁp�qރ_b��}�]mȅ�B�YB����㄁��;̓��2����b�ԙ幦
����ie��0�S֪1�&>�(CM�u>�9��ѶG�Ȱ��,��&�� b�ól��R��\����PH��,ohyӣ��@��M�����U�ĉ��T; c0�:�i��L�"�9iݮb�<���1"��i\"M?x�B\�'f����^�5�������E:}W��)1�˻C�D�O���6؁H"Y�&��"`>_H	FD���%��N������u�����]RyK�x�W���l��"5��3��|��pJ�6��4A��/#���u#Dfe�)�Gh�ɫ���j�0�$n���ƺ�aM]s����B�f��Ǜ�8�5uq���e�z��J�Ci���'�����f�W�n1���M�;�k].�@p���Dɧ�b��$^�?���H����z��'����'�B�G����p�\ZޱT�Ky�p���Q�Z�ׂ�V��M��s�ٗP�5��D4��}Ɵ31|�R��QF�n187�IN�Z�(0��� `�(�
�Hh�GY@9��X,��t�1	B���RRՃ��DNEP7n�B�眃k���G ���o6�.��rdr�Ѐ�绿C�5��0E��X��-	1�Ϯ�YI�����"����%�*�s�Is�f���a�����K�Y�dBF!��H�w<?�`�$'0�4���lda�Ͷ��� ^,V"�Nҿ�wx���0~��Q���S���z�`?!R�����Z%&��Y��F�������m�Vx7�D�)l��� ��L\�NT�go$E�3��x'>HIen��q�)s��u�!�A�X��ʷ�%�>r��l��;	Ra�xO�T[�nٻȘM|�%7>�
��ᗤ�M�9	#��:2d�X�d��� =���Z�߁~��v�ά��Wp�?�G�^��9y��P�NP0�E����5FY칚sS���(h.wmvU�4C�ޞT� ��U�#5氢ЎYg�l�Ǔ,9p��N�r�}�fPz��^��}��[��d�֓i�@��bקُm�vVS\C����L��7�߬���Q�v�"�߁�=�י!�=	6wLTp�)<��:Q픭4�%�㷱\/��[]��Ze�dc�7�X]� ��3�
��H}�o���.w@
���׿ρ@x��y͑T�X| E"�k��x{�?�rE��+��9�ۄ�|��U�u������W⪲�q�r�O`�AA]K�~мi*![�qi(@D��h�ݝ�v�e�;�v'����1cH�7���vr�r���v�G4�D��i����]�G$�Ǭ��Wғ���{��kh�1	�p�9�07o�����4]��tjH�3��H����e2��]�rc�lW��&�Ն���N�kF�
~Ϫ���FC�*IQ| �Wl�s���gB�i��3x�1���-,��@Fx�?�(�q".��f�7�d��2q��m�T�q#D�o���5!��&н�?A�v,��0θ"юrO��e	}�¤Q����4Kž�n)T�����x��8`Ԁ�2�?�I�"Ӓ�n��5�3V�?�P�=XF�Ӝ���Q�O�Ȉk����`c;�B��w���~�?�� �f�\�E<�kL}�s�_��N�?CY���C?؛FeR��B��r�+V�6-�q*2��T�&\�7���>Q:��	|�1.V�Wj-�����쓧�����{��@�=�Y��$A���T�/.��˪f� ��Ic�X�Vz�J3��!�sg�K~�]�j�W�mb���m� P�#�}
��/h�A�4A���c7H�*��#��B+n� `�ʆ$Qu����PN�l<"�|�j!J����o��w���5?9��͐��re	�@=��n��񬐫�5
Ü���l�N��� ���jϤf�&��rwnl�#G�FO�ßBT��})E"�ް"\Jr9���%GF*v�����3EQ���fϕ}�������xr�8��s��{"��h�Q�9�y>�4Z��n]9��'�gc���`�q>��#H�i�ǒR~�4]�Z%�$�w�9�5^(����	Ʋ{j�Lk>*9z��p4����a`s�f`�[������JU���@y� ���鄸���������Z���^����������`�;\e��W�x�p0��(�Y��DX@��?u���?�D�6�ZSA$��� ]�m�	������=M?�v�,L�&��%�o�<)γȟ���&Tǻ2�ť�������e�r%S�=fFmЩ�ql �e�����{d�b��� �/�7Q�P���`\���0�F��Et��
���3_Y�]�� z��=��M�ϟ.$���D��9$� �И��dT������P�L �B�)��Sw����a�����T��ڟ��H�R�e��~��+"�{��5tP�|��RqXrs�xt�N�ņ�/�`}�p���8�WT��-�H١��s(�:c��;n[�+��!��#�@�(�VA�}�����Z�n��7��,��:���?���S���#)L�H�w��t�{�t�M�甂�?>�l��R����I���th�vWCX$�&�mk�'0��E#�����8���ő�t�Ǩ��?��V#H��V�����:�3W�fW �$,G��gLa�L��Ti'}v�8�G����Nx~ìW5X'&t{i.��5�Uy��:����}<�0е�-�wW�c�+E�y���,''xc��	~>�������啴��DDuDm6uӥ�l6�;�9����'7z.�GMB�Ѿ��[kWN��;��f��Ūޙ���M��wT?C�|ħ)�)��ў�J�5�?a&�^8�!��)�z�l�,�������"&3�(�3G9�V���F���e��~�`>|�:��}&L/Y5���lD���˥u��TTręl5�wNIn����8�֕\��	'+{������%�
�� 9! �����I�����Wl�V�Q��΀s"����>�#$}\�1�E5bd�O&B��o���������,&�/f%�U��-�T`2º�e���3H#�r�GP�tsl�T�܌��2CG�B��_����[[�6�5�����(�_�n.g���^i4�$`�G$�ܿߢ	?�*�C��ap�_,�vurN�՛��oN.8>�����9����)�yk����e�_�9"�-�������%嫧#U+מ�.�0�K����<�ʭ���p��r�?D�U����kֺ`ǉS���'�`l�����?h�e��ůt	��[!�^SQo��1�wo�x�a��H�L]���>⾺�,8�$Z�%z-	�XK��N�&�w]��>��'�ٔ)�f|��9��n���kW�F�)a,�`�9�x��%���ܹ�qV�!Ŧ��������Sb��,�q"���� �,l��� �!oI�G&��;j��kQ�������_ʥ������f�JJG ���2RQ���>�Q6e?5�}�;#w���-�V��	�F���4&���L(!{W�{�{�;tJ.�da� �K���	X�\E�#ja�_��T5%v�"�?LE�Nq��505�l��a	���6[Qr8�L����ɀ�&[Nk�j�ၭ��S�VN�EW	dX}3�@�)E�])]o��X)�3ܝ�A�<R����?���]"'H/P���w���^'�d�����P��[Gg�|�@�'1z\K�i#��Ե��ڸ3j-�HWns�N8
�pD kc�����n ������e򵉓Z�q��}Z�<���6�k�C�V8T���a��>H�^p� �%_*��ׯPǧ<A+Lٺӕ�31*�D��Q8�l�`���8=Ϋ�P��n���Gz@�s)X�>yG}�S+�h�L��j�x���������P����Ϳ��S��qr��N�6"I�����%@������L ���|"�f�zg���8n�_a��ˁc��/���xw��璱��p1�TQ�'�ƤĩM���LˢeUd�d}��1��dǖWNn��+��[ˁ^����ѵ��#�^fC��͙��II�⁡��l��������W�28E������{�"0>�;�Ej�L7�S�7Ix�l��]6t1���T��Q1����I�y���}� �E��[$=����Xe�鑏�S�A�ӆ�	�1�%��+��D��J$A��#�¼�&���"���A*;l/T�l�K�1s�&��	��E�Θ�נF��kV�\k�i�#�J�E�؂vmĘ��.�Vw�P�Դ�Hp*����̢ɀ�-K�!K���-xY<QJ��q�-��@�z�������~=6+��kU+�o�)Ν�����
�!;�/��+L��&�j�ڝE��nW���B�)����%�`�;�jq���WE��Ӵ�D��E��ؙQS�L2�O�Cn~��)'�&v�&* �a����`ܱ8�	� ��*��	*����&U�fXċ�|�p�C���	�;~�ȩ@�-<0�*tO_�x.���2��[Lɠ�����<��?^'	��c~ܝ{N�W��*�|>e^��¿�4&0F��VoQ4����2�9V@�٬y_3T�CL����\�����n���x*F�Qn����-�5���sv�@�*���OD�I8��1�U�9Ʃ�D� ���Z�\�	�3���%��.��ƼV�ǩ�sY6���a�;&}v���-�\FעȺa�I�+n�əfX���6S��ǟ5��<����Xn���h��"t~=�F�15��5�al\��wɤ50>���mk4�־M�`�����	&z*�;�{'�{�c�݋��RA�������s�Q �܇!����t�IY3Y;��2+7,[W�UH����c�c�������*�lxIʭ�����w��&t>&�Yi2���A����(r'{���?���$���B9;�Ν*����ņ	�?���^͢f�Q�x(��V�Bo��>��:����	ddIX\A�o@��?�%|;}�L�+�H����E�Khqc~jLd)8�9@�<u�B�_�(��Τ��,��pN��ܩ6`K�m�Ex�ٟ̓y��b�f�5䷱�8���L3�c�j5��� ��P��|�Ϡ�ת	��������N<G�����)�_PT2Ϧ���;b 0uu�\�3���&��8����=AD�Z,��c�ym�7Q�Щ�^z������F�Q��D��pɌQj���p��`u� �L酖q!��[�Z���ࡺ%E�s�Z���h�)b�e�dR�6ʜF@�:J��C���*�_^��&��%g���):H�:x��^�#��Z{�$��5�{�M��|�z�ףC��s��<d�������6q�dS���\���,9AO�kְoRz\�\�x3fy����rHA�ѯ1y��X���
�I{��/�l�f��<h+�LP8��'r�^,D2��r:i�E"���2���n�E$`��4����Mcג�yy�c0��|��sը�oB�����y��_yS�B�>�Ԇ7>5�I����ES ��CVh�1 ��Jml�&�7cY3(<����[���!����.��Cb��Y/f����{z��h?���SϮ!�#~j��L-�~u��9�Þ��ų�sZ�ڊ��h"WݸW9��<!dq�������]
�ݺ��3������C�:�v9���=/��F铓�K��h����m�ݵׇ��:�uǟ58��ɩ�\n@�)d���>�q��|=|���d{�"Yz�j���d��7S>�xX[�8�����E���J����I괅
�?�PY�S���I�AP�ӈ�9�
���ߧeO���Y
�,5:w��/D�����e��@;��V���!mq}���!k{#�V�FB���F͉�Qi:�;'��dv�-��GT���`y�vm��� P���=�U�L5=A<���[�8��i�r�0�đjp£�5��^�ĺ晥�͂I�CJ5wf�*a^�ۤ��Y�a!V�/+�CDw�(\Z�{ݸ`%��?�S��8���B�$s�\�	����h!ZAG�s*�ĩ� �B"��b�=�>H���N@Z�oxk�8CC����'_�m��-�hU���p�z��_gL�#}��_I6��ːX���@V�.uw��0P=�S�Uvg���B�|�wC������a��C��u�U��XfC��=tj��;QesG�Ϥ�Av��U�{��j���M��'�6���W��;^��V����S~h��s�f�_&�����$T��B�q�Mj'�$3a��D���.{���m��.G'r2�rFtB��攢t}�\D[����eAD5����L��:���_G�Gǝ�mw�z<n��|��:s֒���7}Xa"%h彮ʒ������'��@��̠�m���mBC.�y�Z�@��Đ3�^X��&Ns,�4����LAh֕4I������d1Ϭ�ĜWhN[���x~ڥ���d+<l?`d��aF��饌�-�VZAڳ�(�����~X�1H����]>���N�3c��k���-�/G+�N"(pl�G�ٛ.?$�ނ�/5�����)��E�=��u��?�
����ǀfd0C��e�RSd�&�Qݢ��<��UCi]�|��*�S�Z߰�z9D��������S��Fv�T��`�81mغ����{�]C��$���/���	��$��P'�i��72�s�^�&�&j6���p�j��Z�M�IЂ��}��Vi˵�n_xm�'��[�,W�djd�"�A�XZ>��%�K	J���ڞ�	P�Nz�4ct父��$^��`���a�G�#�m#% �lN�`c�.�FD�w�@����K�O���\�G�\!���nA+t��#׏�oX�y��!��>�`���xM��[K5p?���h]{ka�>�ߨ���;����!�'�v/��^���y��#�X�,u�L�|-k� ���t�)����R�%
%t�^�#f�п��-��vw�7z��d-}G�|��F�E��� Gτ�@Ÿ����I�{"�t��t��P��y����H�����]īw��J�e�!���'��!qBy�F%EAea��#֛cd���7��S�
�yY����C�Q̌���F���C*R�\��{��l�Ί�]���Kn�(�˦Ns̈����u���_�S�OoUN��E�,�`Z9D��Q�ek�aϟ(c�Wğ%�z���0A�A]�ƞ!��k���S7��,��<�:��q�"���C��5o�w��f<���27�����eJ�k�i�np���Ǻ!���4��%��v�H���iB�[e2������!��b�5udn|�)񇳹��r�y�ö��D�S[�uE�@M�BGu�i/����hS5�KO�:�d�i�;��7�p��_�s��v܇?����\���U�q���	"���X���)�޳*�)��$�k�{��p�j��� !d9�c:i��a}��e�F�������w��n��_���ExK���������?��`\#~'��V~ ��V��$1�/ +�i>����onM�BR���j�g����I��r����:M�����V�U&�fUx<Fc���P�Մ^�ޤ~�jl���7��l.�Ln�l�ؚ-a�Q�'\Be�M�*o�@H��[8h1��q��ױEӽ��p��|���hn�'A*G�w��2	:�`�/lX�9�p-�U<;
|q��"����d����*��=��{�o�i8�'o�G�ԏ1�x��kb�|�����Q(�l�+��Y��t��UH���y�\�K��e�9�h���F�T�4���w'[���L�:��
,,�р���_���7#zC�d��C=���Pp/1��������ٸ�_����N ���5`,�uKݏ�a�����ը��*�a�$���)�Ջ�8���g������jm:���v�Z���S���H�F�Ȟ��7���;��O���^��()۴���5up��F�����,�:��ΘX�:Cay���!?�=�e�vDX���ȟ�d hs�r�7����/ `�j.������j
���7h�BjD���v��@2꡹����O$1õ=�8:�! %.���s:_G^�����;o]��w����1�|��z��@��v�U���m�1
?��`��< ,����b ���W N'� ��Z��޼B0c��Ae
q�s&gY����H�`�5f�"댫*+�	H^�9�(��:���C&���$Q����]v/%��E�6�k$����x��6��m�*��ʞh�R\��,�
Xn���]*����K����Z���Ӵ�w��t͗����$B:�$�NΊTA�2���*��*��ҥ3֏�.����1�|n�]m]GX�ϐ����I�쩲��%9ֳsE����፮�}�#*V��sg���:&�'C�/G"1��ó,��-� k E� ͷ���by�h�qS�蜏\ǥD���;��s�D��� ��E��L�~���:�70e5
���cY>ҩn�"\���SN <P⍗y=4}�tF�:��d��D�N�v���_:�D��J'�^�;�;֠}�W�+���y������������}r9�_+���X ��B6�,�_]�2���gҜb����`+��6W�L�SjE�v7���#:s�����d`���1���(r}A�����x_
�⣤��ca��a)��3����ـo�Y�R�̨e��Qe}����6�ï�]"amx�AY��<�����xru�i<
39y���%v�r�G�W!�a�K��)����쯿�cNFvc5w��G>߷����Ɨ�زGp�6M��OH�*Y)\���z�#�t8�P��\!�9�E�Q�}��y8�pgnSPM�yED�U��A ��u)�W̨��G�;Gx�>�ׅ�co���Cw+��;N-�uq!��@�o�~Q� ٖ	���`��#��^N�����P�s�B�~�h1�i�2bW�P�1�5�_��≈g�j����A��%tUu�%�m��W�C��I,sB_�_9vY2M7ó�ަ��V����Y�<����?����¶n��K�ޥ�;��q�|����VK�U��X^���&�y��??p��;b���O�zj���"��_�n)ɋ������pt�?���Js�FӖ�&�F��;���b��;�E�΁��OD�*�6iK�V;��Y~{����)��a{7P�"I����c��d������G��J'0�.t?����u�����i��O�L�z.�f#L���bv�v�j�r-z�w�WO5o h&���1�]�r�n�2`7�T^�W'KF�!Y��y�#�8��)\bنC�ff��
��8���۰ȉg�Y�c�9���U+4���u*I%�����#��)
E���3|�.ӣ�(�!�P��z��NL�a����A�J�}���q�=�0�c�]᪼ʽ�ì;h�ra�b�h1���M8�������=	yL���O]�����K �a��.'����T;�T_�C\5����z�;;+%���%pv���|r�2����L��7����f����_���ݥq:��@T�&� �}�[��M���r�'D��B�]��{��"8�H>D���;4�1��?�K� &ɋ��y�)�y��FT.�!�*�*�7Lb0���=h�円�f�}	_��&Y|<�~I��̪E�j~ټ�n,�����!����59�z]�<�d�GI+���� ]4���R���7��{�L�z�)t��1/]��|��g9���.�J^��|�B�6��lK��Z�Q�Kr ����3E1:R���
�Zm�P��	��DB;�^��K�s��7wS|��v�b<�y���`��^��	Ά�F:��޽7�[>������ֈ�|��s�UƜ�3Uەv���fd���r�7�F���K��/�1Ǐw��
z���-�{$�&R��y&R�Sei�9Y�Rr#lr�������64���4	޵%���$.�1�2�tG�UX,�����8@c�\TVZDl�û�1_�'d���^��cp�=ɋ� �J����7�a��(Au�_����E�(�~��r{ L��j�a8N�0�N*��EZ�#�[3ۗ��(BG���"Sa���,�R)��	�"ܢ�øHײ@�U�B��꒯����zFR>Y?#UO
BV8�:wV���VM���2jIs��2�G\�ga_�{U��ՄP�O.��$�L�"���n�e�/b��bp�{5�h�c��߽<ƶ��-ʄ��[��G����bY��,+��-�)��?a:��D�-�e1e�ɻ^N��	
�#'�Bx�')�+"i��c2��aɧ��wu�SE�+�{���!A�Й?��U@��Y:��FA���Y��'�,���w�@�Zև5�ߠ:B��m��?I��/`������?�8����K�ܖ��2�:*��.i����WW��I�1ƒ!4��b���GiL�J^����(�.����T2U���(�%fyxI�[!C��Y�-���s�7�j��Ŀ}�UF�%�,�C���Er��s!�{�0h�[��i�W���-NV;	?��O����  ȼo{�}yN��0r<�M�x[������p§�x��j��#RG+�D�� ������*_Ն��A{����F� T�ïg0�RW��7�%+���}�G�Բ�b/��3Ҧ���/<{���� �V���%7��Ħ(�Y�o����DԗT���>�YF˗ϭ��C#`B�p�-��\��n>�o�ǖ}���Qo`�lG-mQpL�hf�&�lc���r���Y��V}!�I�y�ꛘ�p7Z�H̉Q[2�e<x��E�&���M���0/�#���?Ԗ赉�W���5���#@�E��N�C��W�T:(��$�5�5�w���P����Fj�p�(VF/�+�C�/z%1�B��=��3$$�3�c|�E*�J1m���=��:�X]�j�z�k3��RЋ4�o6��4�Kr�Su�2f�^��4�����\L�/X/���T@H�%��x�n�x�MT#����D��6��{�2s���$���� d�p�!S��z�v�o�����t��n�N�~�mɖ��"� �,p����G��f\��@�L���۽\�#؞E}���c�����6o� ����qR����^�?.��y�a,Fܰe��_P��Q�\O�ꚭ�!@@��Y���8��S?�%Wy�����Cy�TTq�[�,��d�r�$�̊��x1�	�:r#�"�3f�V����t�p�R�e�q� {�T��w���,��2���.<,8^寚��\��Z�x�����Bۑ�]�q�'.;��ߤB��%J��q�Bh�~d�eJ����RC]G%W�}��Zl�pT_w�6s1��d:��`<�ݭ<N13�n�I�����˪��w�p�(�ՕۀI��8�ݓ�a�����3��K8�h���,��>"��|
� Ũ��<�����s'�K
	�ǎ������I�*s���6��V$�l��L��͓7��1n�b�=��->���Lr�4�Լ<���*����� O5�;���5Hl�H\�*0O�f0�鲳�V�3����{.�.C�J��<�	��K��l�	����o�3v���#١x��CU�Q��I�R�|���K6u�e�~�K��fK�F�+�I`�!����;��ͽb5=�$^RВ�g�0X�m�6{���T|��Qn��90��B����Qߦ��V�	B��L9�V�,�4��g~&^s�բ�}Yj�Q�1��`�����X����dgoy0�~j{L��fj���Ô)P+շ��P*y!�w��ԏқb�Vs���
��=D�hcE�5�ѕ0
$9/����@ѽ�y����pE�6'�t,�?'�9) L2�h��p�����ծ�������=�!A) ��
hf�T������ՒU����%�i	= g�������8��$6A���V����7����Ն��*��^���ؼ}�;��|��Q"�㥻.hڸ�N�^'e�|p/g0]gX�rۙ����δ7��N��4;�M�t�(j��_%'8U��E�Ta!l�`Ia��x4|-�K��𼯀�á�x�zt����d`��n����~wv�YMПKd�����L�H�����ȉ�2��0.
��O��x��#������&.r�u80����������s�t��)g�Po((h�5�Ɏ�c�*���:Q_����onϤ��-�Q�H�ݵ4=�2�_�{�c ������B��i�e¹��v�2�:�x�iAGJpQ�M_��4+nO�8t8���C��ϱ�u*��EY��x_V�{m�X@eɯ���ǈm�8�C�����m����������{�+���*�7KZ.���!&-x����"���/�-�b��]$�>�fF���1W�=�s��`?!V�����BA��P����|�ӆ8�~���/2O`ae���z���Tg�z���|�>����ji�q)�q�^']�+�0�����Z�mv�4���r�G"=,'�7�d�,B���sxա�X��O�!p:�lP��X�_7jſ�Q5K�F�+��A�C@���W��<-ɷ���w���֖`A�C�t�p��7�Um>�%��_*g�̸��怂K�c3�[Yy����_;5�ˉ��ysc����a�\R���-�o+�jϧGb��k�K����5:�`����G'�N��Tw�D�`�6rϒ�����Gt{+�l���>��hܲImF!i�;R�C���@+���3@�.X�����D�PD��uQDZ��X���)�8��l���P�-^����'�䕈m���*F��Lq�<8���l��c�ʾ۸�EZ���y2�XJϝ�����\$�֧�A�!>�����^��8f�������u����;��{����&pNH;E�)FXp�iڔi�����{�WJ�gx/��;�띇���'7�cS]�P���Դ>�;�y���ɥ�\�Zc��'��DP�F�X����ֵ�Oc�-�K)�dzz{2R�l��y ��.��,H8h�ݫ)��ŷ{@��wq`S��B�;����3J����A�����&�k�4�9?�W?9�h|��� 냕y�<\fX4��^sj���^8%_\<�*�z��(�9iD�,�-�$(}����%�6]��w$a�������n
�ѱ:A�Jy�� 	��lN�7�,^�����\c�%�Ah��V��Ma� �DsL�9w��"d�逧��\2n�%MO�Q�4�][����ա�����@6���~;�!��WOL���������X܉|�&�o&b��u�TPF���B�A�'������t���ܦŸ�s�)eD�"ڈYG.!<(+��1�wրp��K_
nZ�8to��++s��S�%]���&�~&b�'�:~[�J�ˠJ��� Vmc7]�Q�i��x�\��Fe=�|��ݞ�S��QgI}��mH�D���$¶�n��d^��<��z:R������4�H2a�@q��&p�\A�z8�:Q��/��/}�@jC�<#��!������ohA
���"S� ���`�������>5=E���yݘ"X�葍X���~[�?��p�"�������M��B�;
)Z�Gȵ�r�A���*v�r�c �~�o�WL8���N��1	�ȤVn�p��̓?lw�����rh�d��^z�I��/�|=�`,��	�FSBT�}�Ųj�NY�A��`H�\�	���$`B, �Y�7�5J�̆bAc���͚���r�5��9!���
,�	��� ��*�'��O��Z/ B
I�t�|��lP(����f�%�g�E��6���l�W;�JD�q�:���R����[AT�D_�wzB��D�ܮ���3ڭ2����W�f�F!7�\�#B5+���?I��OYf�)�}Ƨ�~�F?��-���F@oU;`��q�s�A�.�f��δ����3�w�<��^L�Ɍ>r�''�1�>Zkd���V�w�J�z�MA�V��ol�BYﱺ�i:��t�i�;�So�~h�/o�`�ĵ���D|@�"�{�*A�P�+��-`�ٻ��t�k�"������(ַ��^Kh�HS��,rPW�?ߔf�Z�k<<2����~S�b2�'s�8s,uH�V!\��9���́��b�oPo$�_�ū(e<ܒ)��m^N�p�KL_�)��# +��t`}�!�9�;�e!ԡrtI�{�n�8�[�i�Ӊ!��ā�jO�"�B^��ȴ���P,�R�M46^��r4�:�r���M�1�-��7b^N�=�Q��j���׀�����S�����<l�e�h"%=�%4������O����u"��e2�k&����\��~\��I|�l'-���g�����)�Uh/�_s�a�
Z���������:$��AB��V&c�3G3�=��_����r������9F��XowTXg�M3i���p��ק��xK�����n��-m�6i�%��g,`v@�5S1��0�m��A_�.~сh[�t����Jx�=��x܋0m�Ä���%��%��4v��u��X\��S��0j���yեu���t�0�m�E���o±)���&��fN'�O��F�J&�&�6�G��%)6T�S�ipS����`�yz���I��J2no���Q?�$除���w�����щ��⩺�����ې��y�[�"�3���K�Џ�D0�)�2G�+���(���c���Z׎1@��;�� 튔�G�=/��OE�H���T�r>��RT=�T���5{�EF��x�v
f�wώ�u6R+s!W����lU]�ygV�iX�4�c��,1�Z�iz�Q�㋊.���p\%���� Ȍ�2�����6�7�^_qH��_����U���H4{���(�52Ѩ��2��f���S��sxڶ�E��rI4��_�$�7WE�Ng�{+�+�W�S��TP�	\�KJ˸��4���W:�Xf{D	��s�hN:�}¾�����睂�!��2�}#0���]�,�>t�2�����3Q��?��>]�y��]�,���'��/6����VXƧϒ��A����ν���E�9.cf(��󦗄��V���4xs�?����7VrV�{��ƅ�������@i��`��]:�5��U��>���]+I��4�F��ǐ��Y��4e�}G�!�Ԏ�՗�8^|�峹�m�eP��L����W2�� �=6�Ž�q �(�1�%�lmb��'b:�s3��h�Oe��B�3uAY��}[ј��/�����e���~MI,���R��%�����)T��S�4�������pJ��9S�AN��;?�-;�e@�Ʌ�Ç��{�yl��δ��8���Z�䀂Н�A"��K�"������Q H�16�ޡ,1%�%�k�uoԫW�W(���<��4�<�â��>������֍Pc	p��y��29{}�z���M�ZEy�z;@i�����3�n�@R}gsk��.i� ���$se��Y�����>�Բ�?�^lX�5u����Tg����G�<��������Gݍ+?mqw*����`$�� -� !к�I�hZ�#����p6�߈�U�Z+�_m���f,�18�l���u�H�k�R�c���������	������d�6�"K�R��T�&�py_]�;H����~Fg{d���uA�M�e��y�[�@�gQ��� �,3|5�S-g�]�UA��|q�~E�+ּ�\�!Z}�S�~IE���L�{���U^Ӿ�4n���iJ�s�݋��ֻ�oO��7E��q����Y�`�$�4t�o�c<D����f}���a��-P���N�����%�;Ѳ�[�8�(Q�u�6:cT�Y�^t���eDvv0D$~H���
�m�o�YtcP�p�����:�s�r��-g
=T����-r
��(g�/d�Z�+$���`��jGX=Cu%�p��*dpg�,�kE�	)�;W���+��(_#!�s�d3�u��(��f�����Y2�=ĕ��~P?����P����ӹ�x�K���O��	M-g�Q�;:�	�=� ���@U�ޠ�C��t�Ҧ�x�܂�R�c _Ii�ĵt��7E���At�@�Mg��FF�x1)s��ΘF�l����G�7�F<׭���/]�̓BS�ͬ�/�[�BA1b0{�kU&�3PJj�(�C^�x1�2���i
g���+<P�>���V��� #��_/���*��$��<���w��=������3W�bgi�Ƈ|����R˶[�A��H���"3z�ȴ�Y�=D�'m"|��L�� `D�z7i�c����h�o��vHQ���`<8+t��7Pi 3�����_�|���n4'���������io#H$�����e�>�A��P�uO8M� �j�㻯R�����g�X�4^Z��"f��f~��~�d66Z/l��/RݗXո_��8�w�/x���)�Վ<�����F�8�;��7�%����������
�m�v/Ԑ?��ٵ����PmG�c�C��<&{�\��B��X��I�5ۏ�p��̄!l��7��$N$��[K�%����v�˩�/��xlͪ{n]�W�u
�3�i�KX�ѷ�7&��V�J =��+x��*����"b�1��N�qU��o�'�,�ʐ�d{]���>}́YPN�!l�T�� OI��B"�\�;��lnз$�|��X��鲔m�1��Ѫ�����͹�V�T�.��b��xIZ<e���I"��	����<�����<�6:bh�&b�*��s$�(�.hg�|���Fk3<��~�Y�'�;�y����2�&�м�����$�����2��weFƣ9�����LHK;���ZbG��-��V�}�t��N~/돧��؎%��UH���U�il+��{��`�g��,R��G�g�ևl�Ёy^�3zB�e�|9��%��)Q�>�6S$��O�q�	�@���I����JC��V8�
C���&�>bօ!�G�&��a���$:�G�,"X�?ƺ(?Σ�>^$t��m���b�$·��qg��G��g&t�L�敃��%�	z�s����{�o_v�RԔ}�~^3[��SQ�Qd�w���(]����&�n"�ͼ�40�JɡBu| 8M����&Ҳ�0�Z�r�Hˋ�W ���@#�:c�^2+��š�g�����$�4ѡ��4��k�7W���- �0#]0���m��0�Q�.�%�����ā�2d�G�	��+F�!U�rl���|�(`Q���h�����������_xHִ�$Z�_1��`�쀮P�\6b��ҿ�����>4�]���]�v9gC䮌��U�	E���<`��Bqt���	[�R��������� �}�װVl�F��n>G�
��j �W�n��+�k����!���p����~L��ߒF���x�.u�j�(��o}�d��`#7Eeb�:줄� �$�4fz+������y�:cM�j�DS黨l���W#��O�{y��ڜW�joMn_
�>È{,0p�&�z.w+��{�s��³�.��@��q!�Z0�$��?.ģ���0ʯN\���S0�w>Nz���v�q)KmD�tab�A4W�G�F->�1��
�2��
����'t3I�e&b���-�b�)���6QZ{��]��e��e7V\n���C:��7�>?y���e);��o�� ĭaA<�4�.޹ɵ�%Z�\��	y�Kv)�k�,�߻��77��� �$��2%
d��Q��Q��n�NGrV�}'�x�7�l����_H���F_K$�˵h�gx��c��%{��l̻^��=��ꀤl�Pq�tMhO�J
g��B��ې�6�%�T�$q�3uʹi_��e������u2JV�-QB�U�`z�$W��]2I>��2U��.���o��,c#Y�1yj2�ꎕ#��г���r�_ �'pGh�x㚅�W���V��qf��*6��W������k7���m>_4p9���핫��~ac��r�� l��49�V�6㟁�@`�d�p��=�*Y5)UXd���%��>������<��[� �jP���&�t�:��!"@����]	��k<|�7����ĉR��f+�i�yEz;�j	K#�E�T�L�}�-�x ���~-G�l��(��s,��l���1��>�E�l�h�F[
�	 >@�q5!�D�F��(��E�E�������1�.GA�?%��(ԙ���W=tf P��g2�X����˓����@o��$e�*(����!B�gȪ�	��ʄ.�|IU��4)���@��JȜ=��!b�k�D��hf*"��]�P�X��(QM��t��}ݑ���^�?�C��2"GͰr����!M�T�}��8G!�3 �:얫L���sU)�A
 �ؗ�~.:�|	���MQV�_�X��9��O=V���_f� *�1[1wkEU ��5tf0S?�E�����X�]���m�m��|?�K�`04}�~M}���t/4��h(M���G�썵Gc%[�Y�`Y��(Q�T��fQ��fhWRU~���==�DT�[6BYG�C�N�q]�e��������-i��AM����v��MHY�>�h`�l�3X8�3��Yn5�����>:��GR�'lkv�����<h�]M�N��Aɒ��^����6�v�2C����
2�N�4ʏ���$�غT�k>p��$�_l��c�n�Vo�eSC����ﺍ�x�mޤ38�ZG�'��l���>(��|Ήך�]!�LQs �H�I���`�t�|SK�Ɠ�1�W3��^8�%'L��i�Ʉ zm+�ƻ������^���/�ZV��Su�]G-�5��A�Bav�ҕ��F)8�μ��9�"IɃ�QԀi4@DA���C��~\�*Ne�9ʷ�w��_<7��W�\	���xTQ���n�@k|��&�x�q��H�C2 m_�U�αX�v�(�{ԃ�	�Fj��|���		�Tȸ�x������IT��rJ��� �k/4Y�7��B��G��8�9b.�n�Ȯם�*i��&�ܪdi�t7EcB&oX2�Z�&�&�O�����:aW��w�w�̊26l=���vgKl�L���O�J���E�G�C��*B��3g"��Q��3����,F&�J0����gȞ�ֽ�,��N8Drhr,;��n�R>�v�Ž��"Q[���:���S�$��A�7�I�ho�g�QV�?>C��VJ�|8`�np�$�pN΂��ԅ7gF���EM����3햀v��{%�͗WA���v����3��G'F��D1�Š�+R��p�$/uc�k���YL��,�g�����㏯�t��t����<������|w�����'Ua�ڹ�՚�l��jX@��8��Ag�N춂B&@�@���-m;xx:�3VT�2����Lq���&Op�k�ŷ��s�Sl��ϱ@�W���`
J���d��,�RZ~gfa:���N3��0DR7r�����& ��
C/l�:)����Vd�� C( L!Ѱ!k��p��0��B��}���x���~����ښ0})�'���E^z���D��͞$ڽr��q�o�u���C���(@�3*{�.&��M���Y�ĭd�䴢�w�W�
6_��f��d�M�R����>��ΊΦ��<}��a�U�=�E�+j� Ե�C5�-����=W��W\�6���X��<C>9��D�tծ���'֒	�r
|U��|b �s�����W�ե0C,;5������V�h�H��J��Q5r���s��*���%�%.����CU,m���[E4�1/���G��[����W=�R9�����E�Tc�V	��\k��4�^�}�g�#���$?�N� �*���d�>����^,��D�����H�+��"C�h�{@�ia���K6�\Ƞ��ꣷ��l�yP�n0rtt-]Å_��fġ,�WbQ;G�6)F,f˃���YJ������yn����2f^jP��L�pN\
!N�_��04������قJ�L��p��eS�lq���F���0յ�^�����e������w=�$�g��N�80V��@���s�����T��������;(*F�Y�nu��sS,�7S�ɨ
[:��,��v�bF}a��",�K�OF 8濯9���ή������[�f�U̝�k���J5@�Ov�P���M�4�<0����I_�}�	�.��+55���E�g� d�m�`�L��	�oi q��(?��-P��iH#�7��m�~4	���|�`���f"��ܮ������Tp�}��O�"_Lpa�8� 3G�r�n%X8���+H}in��)��|!�!���T��f�=Ԃ�q����8��X&���<Bz9��D�� I����D!�r��2��ۚ4������({8��/���������G��H������O�, B�?�'��+��F�4ɛѶ:����R����/�m��A�,R���=�LL�����j� l�ʁD���W>�1�eΗ<Z�3�F��Sa�_��3�r$jՃ
�����W��dZ�ˆL&��tC���Y���u�_��&ƁT�د��˰o�-W�nS�%At|�)���k�����W�I?B�4?��$">��"���A8;Z3�#�І���G��J�p�{)��"1)�U�ʰ����Cx�8�'ep0���m�h��.$�!�HeJ�˫���r��Wj
H���;�o!�`u���>�r�3���9/e��|W��r&��Ե_+�Ģ�sΎ�x9�5�CU�*S1LS�����g���g��q�r�p}P�Ԩ>���7�<�z?�x/.��'�EM�%@\=-{MYVܺ��k��Dw��j|e٩<�ŀխ9�p5C,4i .N]�<lp�+�L�V�hܘ�*�:8�S��7�="�=��	^����Kk픆y4/�͛���.hq��'_AHۏ��oC a�cd8 ��`^PM��}�s1)m�1a�m������^3({#۠��B�i�Mo��̠!$P��VX��ը2�=]�����x��p�K��P���JW�I�pvQ�nM�K3ut�����׃�R�xܩ 0�:�pg�E�7��lP��(��gl^��J��)qUw�>�6��?�6�@KH��~�U,R�G⴦E�{�C�KW���«O���f�{��~��E�r�BWe����J���i9�s��(�& ��<��gC�jƭ����G�z��l��+)Rif�g��ɰ%Q��'�$sMFsSF��ZB�f2.d��M9ְ[����3�p��m�oX�0���x�U�&�W��V�3kn$fuXX2�fk`4%w��"H�-��:� ��,{;9͠�B�'Z/�
B3� �Ւ�|�t)8^��B�sT}�C��D�C7�AU���#�F?���ƛ�NG�CU됌��NS�ӑ�v��{ܒ m#�
FN�V�����(���dB����W�猙����W0�K솟���~�U?�m�N��]&�f%T:��#�-�;�ɊQ[}���e\I��N.�p�����0�T*���N�F;;Ż��B�fj3Anml	��K�V&�"����qa�C��T��uʧ�j�l�2��vk8`3-7������R,b$������a���PJ+M:�G�}�B* b"Cb��>�L�H�� ��B	=������S�p��a���[�3�W���H��Q�CMC��/|� �1���T���^���D]�]�;���"IDEO�.G��D��H���cP^IN��Y6�A�vN��F���ۥx��#e�B
�G�b�K�5�L_L���qq�x��B����qPn�aÞ�@��/�xVe2W����g�\M �=�
�?��NM�e���� �]��A?l�@>�}���+J��H�����M��4,�k7n�m�V�P������1�A	j��nk�k�T~�W�Q��EJE�Y�#(G���K�D���71�,G�r���6�U��L�
\'�H�ŝ�p:�����ŧ[��m���G%�s���DZz�
t����j����}�M��!�7��@Тҏ������k#DSSi��Ϣ�ܫ���i���Q���=y���Ų�?µ�=kF�%(塈}"I�+Q��qIˉt"?F.�k�pק�4�q�IW9�xp�S��U,��]PX�@�.H��p�7�ؠPx�� 7��w��.oU��ں�ړd�#{�bgn���ʹ�`��A��l���U:�G`�l�i��S=�!њ���ơ�ЏH��ꓠü��϶ˬ &.p�J{���6y4�a8������"{�)#� k<�.5���V� %C���#q���-C��q��m����/��
(��$��.g���ήӬ�:@yr�l��6�t|��o<ٓW�K�Ѻ�������ŵTVFB�	�5T���vI�Ƿ�X�)��9�W���d=�=O��7
"��qG���Dsh�m�]`���廝�)
�Z�xkiI��L��7�2B�#Suǲ�;��A�W9c���όj׼D�y6���}.�(�c��V6�t���~�6�t9]�c����^�Ko��l]-K��ُ`lF':���TC'���34��ܼ
1�_lt2}(y1����$�,��zQ�>����]/�F�8G����`\����l���9�w�NE�����*u��۾}�[�*w����b�3�0P4JƏ9пF)H��������Xv�*�A`àJ�lB-�@�TWi�W�j���$�tX� ��ͣZ�
���C�v�cy[�a� i ����2�ɤ�$��4���(��Z��5�(眱\���~E�୰��]=�`�;�XK�$����T�7v�N��Q&7FbJ1g�x�����rA�|ng�K�5�EoG�O�F�(�0��Ӻ�y"q��{���$�?�8͕ϳϺx�3�� �\��x��9�0�^�H�ɱ���\��ю��*����!�jV�㭻	5��!�թ2٩��6�x<�<23�s��؁��E�z7��%�
1V<��Z�n��?T��	������J�ʙ��x���9M>m&��f}_���	�F7�����w�,ry;��������Pɵ7�	��y:WµshZ�mn�~���i�x7iT{�j#�d�/�~>���v�,�u����]D�4G�l䵚1w0��V3!=y����	1�;R1�n�3�����0��޹�8�}��๣�����h_)q��%�>pxɾ����W��"��9ߤ-D:u��}�/\b�R��bL�S-S��*�+�o����8��^ed+&w`h!s\hE��9Ay(t�>����:�>�JSſ�i���R:W��?K�+v�VCq3�[�c�(WO�N�F{��i=j�M�p����;�4#�b$�G�2f�Uf�$���F���|� ��5�7�:�����~uq�S��Ehjt���*���ARJ��p�QD zR������W�.#Xu��>���0a©l�;Q+��N�Es@M<����a���Gi[,}:�ڶ_��o�cx)h����T�����0��2�t�쨟i�a�X�21�[>-��~����>|]�
�w�:r����d��V+�$̙�����ۋͺo�.&��_�[6�Q�i22���e��m���~���`����E��]�#�J��(����������lf�x����m>�_�6���|���^L	v��P��;��?�!��Z�=7ӓ�v��(M�J��:�d^TN��Q��I�N��o���ח�?�<��b-k���~����4$�\-��V7�b)�@P��$՜�3: �5A7XMS�j=:����7;G�˪�qeWG�>{��zc�3��m��m��%QX�-����A�|���e������~.<��or�^2mx؉Q�w��=��oV�4�����zbV��J��������cU}xhE=Z���V��qE���.�T+oqk������7U,�$r��6 �G<�F'���ː�A5���]o�9�|���fK	T�H�c_ހ�?R�5�]�9`!D(<3�Q9c�x�&SRݼ��W��̼"�J��-��l�Pd�1�J���ܨ�w� 5�ړ��H@B����$�;PF��|ufk��vo��A����B������ 2~"o!c�5Y
@Lc��h��@��k��<e1A�i0\������ۃ�:����%SY�,�N
���P�o,UF��"v�ǅ#0�a��bx�N�n��6������B��t*��&�����14��iX2�A�,�P����7��}#ƀ-��'g��cOŎ'��~l�˂F������N�idI��A�{b�Sm,r!�,4�gC�wr��z�Z��7v�5�E�dh��U���\��mO�ˑ���ۄ��is��jf���g����c(�a�	h80�|I�t[�p;�?zG��[��Ҭ��	���#L	�I�����e������%�	�K2�h��p4h��G�	5���)1������{2E����^*ꃒ�پ��L�2󋂃�~^�^5D�_�j4۴c�&z+u�%rې��n���u�	|j��I
�hȒ�%���TNQ��<�5�(*4�d)��qh�lJ�������^����)�.,j��!�YI��8�%L�h��0z�_��J{��,����0�a�!���gZ@|�&?�m?0��W�խ����|���d�7����؅+d��Y�ـ`u��k)ue��|�9��Ż}�,`Z�5�b�EꇇI�I�G�BڌK�{�Y��_Wt�t��n)d�ɯ��U.~a&gs�Ɋ|���%ȴ=/��E����H� �!F����a�e�a'�����3���٦I�M��B�x��+��X_�=Ɣ��B敠�^=��!�W��R�^r�yP��+�fH|��f�b����k��	Y��b��W�����E��2�:S���a�(���U9�q׼H�,>pNJ�KR"�0�/���Z��FO'�5�a�����ǧ���^G�kO��g��Jڵ���� �������V���-�c�U��t_bZ��L���q�U�
��2�����(���m -��A�=����<����f�sU��p�P�ץ�4r'w�2'���'i�;A�|�����-�I5�#P	��)��t�}�3[�����)��+�{f~��誋�v��+�AO8�9ׇ3c;�Wy�k^����I%ڨZ;s�'��bÑ�8��,8yO�d�X���sTK�#��1SF90E�RG�7�J}8�T����u^.��V�z�G�����1 ¦��"<�ڵ^=$$y�dT2@�`�%�I�-���ҘVGH,�5e�Vs9��I�/��~d��r,��3���'^������Ų��<�h��î.n3؉�r�4#��G3 �EeV7%١�����YX���l�X�["���-����PX���Z%����K�38��8QrK�u���d-$o[��=�4�3�oU��f(4.�Φ���N�
�������n�%���p{h�-�5Q�@��ؓ�5���ݝ,�ʭ�u���IK�b$o0���]��/>lQ�?c�eGRT�S<&�P�珻KҒ���|�7�H&����8DV���ʹYivs�y����I�w���Y%�L��Ӌ!j��0�Q���-SC��F��a�C�Q�	T���ޗԴ�;+4��m��'yl����A��D�������{p�s�U섾�>��Ӡ�[��ZD�����Wlh���趏�.T��j��I{�����eI�V�d���g;��K��6A�(ޭݤ)�04�M7p�<!�����:K���ؿ�KOs<�g�Y��d�K�d�d�mqۅ(�Sak�I�;#�5�
�4��1�L����8G�K�R��/��3ok�)$�l��@c����g�|�!$}\�X���;=R�%��x�aD@��fM�X��9��#V%��bh3!��P���_0�A�%�xβ�v\��H� 0�;��Bi�$Lך��dW<�N�$��ņ�n�jڇP�GU��~�dJ9%/h;���^�9����NO�f� <�T

��跈}���"t�.Mn��8���8~�*Z��Ϲ�abi5�ɾ8�l]z���*r���-� >�}�*�!,{��GT��	�	��-I�l��a}Ʈ�B���E���V3(�dG�l�Q�Ѥ����Mi��|i��$�2{ɋ�k,K�i4� �Y��W�t?��j�7+/w�A��9�	���.)?�m�QE�rԭ�v���/�z��T=g�{�J������Nt����R:���b�1����rd�ˀ*�u��`	�1���c��O떶*���Q��l��ܯ���S���3��3��zB�:�_	L)ҟ(��/��.T�7<D�2�Sv�iZ��}O�s&�4h0+89���]z�Y*�r�WP��8�h�J�>A&��W���)w��5���Em\�r�V@��p��O����gQ��|�t������A	��9���pܭ���g����J�T�c���$�)��E@YU'��ݽXw�*���[k^@�Sޥ���/�9��^��\�W�2�4@��4z��侩dm�D���?�T�\ K-ܛ�@&��0���-\#��
rS��@�F���j����3� ?rL82%�]�85+0c?���YP��o��ː%E�j�ept��Q�`'��_8r���"x�ÓvN����5�²�SW�[X��)��e���c�*�{�j��o�m�����o|r��!�1���[]�:N��"-��[Ā����s)��Safq4i��(u�m���cȘo�-)� U��J��9�h���}[i�0��ԟ�җhV)���i��7x�b��*&C/�:J.�����ig�J�u�yr�$�v�H! ��p)I��	���4k4���!ޑWѕ*Eu^���(ʜ�@��T��Q�6N��ѤӦʢ}�xV�R��T�0�a+������!G�z�� (�{�i"��Ƨz0�J�#�!�T��%H/�����~L�A5��r��+���<	b�LH�._Lk?�vЗ��d�#K�̞��CL�_�Hғ��\�?�,	:!� �aa��l�tx#;�`�<6������+�5�](�uΦ�N�<�]̩�9g�WT�_�'�(�	�p[I�`�� ��2º������9vċ</
N4Et��l��o ]�1�gX?����=��:4Z>۷9��M��D��Ǥej�?Y���'1����"�ǖ3�x4��g�����p���v����&����@�"��(:���(qq+��R�6�'�eJ��NSi�;�����P��x�������{(��2����u�xj�m��`;D-�����V��\X��n�9��ў	�
������@��H~���?�N��y�kw�QA�0��|����P�0%��0܁o���ы~�[~'#�,ɝ�JBG;&�n���ɌpP��Dc_��BĿ/���fZ>���(��:z�˕5�����N��,�C�.��W �}}\�hf����0~���T�5z2�Y�^͏�-����n�ȥ���`����Yv����'_E2:��Uk���7�o:̆KS�v<��j�b����$��41�N~�X����%�� �T��bm`�����B U�d)�m	/���W�򝥃��ߐx*t�FM�۴8G�(�����;� ����y����<U`���*��d�m�xw�N�1e]E(M���M�5oj��{X����������B�pΑ�$�M���E�M�U��ʤ�0�*3N4h����?�ssV�0A�Y�9sHGg|O[��_�ل��	Ω�K���Dʢ�S�
���^��K���O.�ې���3��љSE]�IY������}$�M��g�O[l\�
q����Uk}^.WN�������.|�b��9�\>�S"�i1c��-���,$/^��v�լ����_���n�!<� ���q�e�k!E�Y��ǯ�=ԁ�ߡ/�y���W.�/���d�bF�����h�͐�SZx�N����壶�/�;;�gˈ�éK.�w�b��x��6�W��^b���"4��d�#��F�J���� ɣ@�cB� ٯ�*��	�˧�@qRՒS������(�\��,�T����W�H�,��z��\�!��f�H�A8�"	��D��7����$G��J��UX�M2��tx+<}
,ə�ܗ��2���6�j���r�#��!�;�Bz{i��U�a���pqaZ���0�>���|�޴�3��/ZⱠ�<=����� O�<2mqE�uA�kLei&/�jI�o���չM���=�4���� e���k������oLWvD���X����R�!���`�ӿ�����n)G
4Hrj9�W����V@��a�FB�tb6A�q��A׬-߉:x���饟�Z���|�b����}��~i�΁z���\4��}�d�K��ʼ�U����g����F�{��X]9���<��tj��C��VBK�6�Z2a=�C>���WdW�S��#]65;3���)�֧�i���j�2��}E�[�DA0�q�h<�P��1��$ *z5d҉�_E:!¾S)QJ�h�֙���'e��@f���U�		�U���}n%,E>dZ>-����jq�๲*��q��6WW6�#Q|����=H �|m��7��3Y����d��.�oD���
P��Q��8=�R�
#��@<X�C�v��!����U���}�l�� (����F�ifB�n��p{��Π���\1	_�E6#��mi��9{�Tny�F���pcG�7n���˸�T-��`��i�A#��n�3��s/�qy��m}�� @6���eA����H���3�0�BB�W����/� ��9
֏���?��xO{\Xq���f�F�� ȱ��f�q�E�,��O7tM�`�@�E����.�xxǙW�P:,��ס����cu2�(Q��o�ISЍ���8\V��k���X+n_񭷯�q@E��հ��	�.�vyjEw�ɔV�+ʑ>���XY8�ß��w��x�bw���y�Q���y kh�<[�K�I�Z^¸d�Y���f=] ����)0�k.о�#�(Eh��d������X��mQu�F{�KS�LZ�<#At�̰_��מ��/	�*�E�n����V�_����s�$vL�F� �cW��1��6� ��ݑ�E���VO�a��:G^�]J�n1s|�%�4�v2K�СP#?���r&��=��w��L�B�GO~PQ?+�Jd	��
�s� �?XO،@�����H��Oƅ����Fy������N�JYB��M"C�Ʒ�0�A�
m"���"k�<�͌,uDh�ii�G%t�CF��s[��#��NH����6+a��
���g��1�ŗ�C�E�Y�Ӷe���o4���K��E�{�;�JI�PƇ+�bn��,<�Uz���g�5��Y��^3�����9K=L�*g���
..�9|9h��m�2q��2�f��|��b|��9}h�8�7��#��S�Y���a�|��KWS���G� ��b��A�Z9�y`C���|��3�ۼ���鯇h�ù�"�Ӂ�r�X�5:�L�ɩT�U��<'��$G��?�1��F�OQ�Ih/�/�3�=�Ճ�qP����Գ����'�F�����@E� a����JR��ȕ� ����i���%C��hr��G�]����GW�k< ��tq���� ��?���χdd��
���^k3�K-V�+b�LDd���W9�JT55J�`�����-�L��B�-v�~g�߂�[M�~��N~�aHTw�?�C\��y:�A�8p��p=[��|�q��{�!1ZDڌk]x���sl)%wgU����tGO�����w�|��Fq�3
���	����r����@��?�x0�b���A\�ʞMC��5_u�Qs�����7(+���)�'�1+�|���$������r���/di�bn���ŉS�����Z�_?�����1�^�j��Z�xT�R�i��G1�;��cA"�'1�Ǩ���8v����[x\��6�.mъ2�Ϛ�+�O%��4!���4���-�Ho�z���7�X9),�3@&����0�0;34&��6�((g�'T��f��mf�ߑ�k��Ƭ�-�x  �7�Y��؆�¼#����w�D� e��ZR>��2 *���s�]>�� _�9:��y�c���42�X����7��f� %��(��[Kk%����a���&��Q@RD��
��3�� �ޠ���Q�xW�M�=�QL0�<�2+�5�<WK4GIΜ�Pj��G�,	u�~�o8����kUF#��vQo��5MIo�T_^(P��&�o2Z��m���`��tJ,Z{�o͗�~�L�mqDX��+=b���W��\=M:����X[�-�l���@r}<]� s�N��ǆ�
�Db��(����q�Ep�g @A Źϓ/��	 v��a#b����F����+1n�׿�B6B�g�h&*
�"�J	;������o2w�a�z,_I↪_�B�J� |�έ���h�S፞�����=��X:N�`��e�z~��FȽ�5v�YG��q/�}�����%���E��oK�F²zWj��k|��lY?�:zt��R�N~V��uƯ!utN%�
����)���R>=��ka��:���5��"�y��$���4�C �	F��d�+�����mF�����"v�Z�Ƒ�@@�Q��7���_uM��B�)�s����WH6PZ(C��c����V��0y�k�D�W���!b�'�s>_�q�{�C�DF=M�󃒱o���s�H�È���I���0���mS��v���F�nϜ#���=/j����ʇ�i����向�FH^VTw�K\�UE�9��� 3��#R�%ScA���K�g�@�M�A>_4�m9c��Yi'`0�E�������C���T���,u��Wh���[kTI��8�A��cP^�D/�;9+��Z��tB���>�q� f�&A]�x�Ѕ]U礣���p�����EW3���r��5��"J�т��62]�e�׃M�JII���g"[�a�'�H{�"G������2/�:°�f���"����e���_�D�}ц��D��Щ�!K��I�	����튩�?)g��R�[K�L�>�4���:���M�%�~j!@~�	c���LPSɪ��O�
��(�TD
���(K'�g'\��i\���O 2s���j�k�c���0��捭��Ri���et^���[�đSg�x>��abn{�5��;z�����ؔ1�g �{�0�fm���un_R����{�J
R�F���6��4��>>�[�!�D+Qc� �7����z~�S�:�%g���*����V��m���D�Y2`��u�I���&\����so�(��.�<=]�>
��[J/��8�bJ�����{�Y�v��y?�Rl
�,�.��(0���yf�ӓd�:�H����R5��i=6�9 }^�5�������ߨ�%<����=Q��M�g���/�#��γ�Ha�~J�������W8-i����K����Dw��a������ƒ��}�����Ym�R5A�B�ƹ��8�v�I��V3W:�K���fNz6�󂂹c�����Z!OQR~���K&�;+޸<�=�RD�4�1��&��M5!������f�l����<�������]�'�D�6&8���R�5b-|a9��R-��#O��=�1���I���d1������iVǂd7��T�O�vB�?���%�1�?�:�&6s� Co�E���ːx|��U�R��f>����L�F#��ٛ����	a����2_����Z�|@�j�+������4%{cb���mQ����&������t}|�v�[Q�h��݈��X5�p���d����?��囒�nd�$��.����v��/�8�T�O��P�:J:xs�|PGz���\�+/?�M���YST�&</u&jA���>'G�J�T�a�pa�3�FU$1+ֶ#s�Enr�t%�*�
� l�ϐ�I�y�7e�"�ʲ�4�(�mU�Lg�15g�Ԋ�s�/�zZ@^����0`��5)b�b��6Ue�	[E��X.�s�= �ce��o53m�z�����s��N�����͹�쨋N�uB���PrG!j&�婤��K�[�2�㦕hl�X}�����Y����Yt�O�е*̜��d���@���)�zZ�$+���c�o0O��yߪ�'�'EL�Q:���Q=��G�L!9����q��pe�E��b�0����;̐[dݖ��c6�<���p���k�F��p'�h���l�x*W�j��A��LW_]�Gq��/��2	~a�����n�p�Y�Ă�E�N�J���Ć������mg��I	�W�{�Ȃ	�g�ϗ���G�bp��"�N���I���X��z�O|2�a�ǜ:X��VO̩X���C��JʼG"J��E���vS�M�� M�Y�^�� !t�r�~����YHD�d��4�v�O�R,W\�߹[{���f���f+X���J!$�8�*����H��ݿ��vG(�`4��R�6'������EZ������&<�i���YV�"I[
�w	�Ŝ'�����R�ŗ���������q^���T0fx�>l%S� ��$L�f���j% �g���	b~��,00e����KQ6lw�0E:��Z'�T�q(b�
uP�[�8YtTV\��&���r%���{��E��l�{��o�t���7-��Å	���OcsF����S褪\5�|�L�#V�� �r`ΘPw\����9�t���a�^A���� �C�嘡t�Ks��W���I5CpE���@M�{J�K��|�wE�����<5�$p:Q���s ڐ{��P������I�򦯳=f�c�����W�{���&:�E������GL�?**c�f�� l�n��R �c�M�yu���S\�O�K�����1��-b�N g�Ŝ����<��]H��C��0lT������a��%�̷G�"b~[X�p�\쥚$��(��I�ne	��=�ʭ��-ү�[���k�3N�u�9S���H.$U=��(ؐ�3r������ �����	Gy�|ɘ�`
�udя
e�2 H�rܛ�1�o-��|o���&� �fsS�$<g��5|���
����!�a��u*�}��'���W�!d@.�dj;w�����F"x�o�dO�p��s��¾1؇�4Y���
ΣU_�:L��o���w���&ΰ�U� �L�Q��3e��<x�>8���B��F�՝j����l�%{��q���yJ�,p����Cl
�D��g.hQujL��N0���Ap�����QP.:{�@�x6#u.�)��D���|�dv�jn�ӈ7"�b�)�Y�B��9]��6�p����vߞ�q���+��G�"�:�oc�O�s}�b�	�w�czM�])�ra�gIޮ(5ZT��:-�e�ֆ$����p��x�l��I�e�
�'\kh�=r�����sk��4�� {qp�d*�pU����2J�l>¡�PqL���'`EPٛ��8�:9?����"�܂U7�����{�ֆ�5�s������Ö�6E0g_�r��,�6l�X������k�J}"e�&v��$�y��l%�r$��1ݸy���H�E4���LPi�������Ԟ�RC�t�@+��^BF�Tj����󏻬�9������A�?v/-	$�+��2�c����jbf��q��� �A0L�g(���6b3;���oou��
�ܟ���tu�Zi���-�d��<�ߜ!�g���k &x��>��Np��%��0t牂���pwy=����~7�g>;ݪ)ԄzS��Rh�#���A�οa1�!p�j< �~X�A�	��ܥ���o�q�}�E����[<��`���~��П�Jm��T���?�X"	��wkH�5'����!�۩c *�����	mo�}�Ly|5?��t")9���1��,))���k��D���x�1� �4����7KV�"��b��� ޸��y�A8�����=3h�JYp|����! A�o����]��M$����zVehD>Bt��sW�U�K��щ;������7�m 醄�la�/-�%m�o�p�g�7�c�X�����R�w�<1(̻�l�0��2���4���W���@Z;>�dw�ç8Si��YZ��Ê��N-T	+?S���*�����d(�G�ӈ����B�I��G���+��yXUW=��| u犺j�l�13x�_�o'�(���6��v������+2�L"�ŀ'J��n��?��� ,{�<��u��zq�&PC�o��B�I�7P����]C]W���AM�&:��g�Sp<�.E�?>"n�h��U�3#cZ�4'_e�TOp8+(�HCI���^J�b@k6�iY�*c�4Rz|+�Oi`ChQKg5Y:E,�Re�xF�'Z��q��Q�8��˩��m�$�i\Ψ�u�C�����Y�tc_�٥��h��٠AQ1���~�����`�4����Ȏ"R7�NY=Wt"��^.�x�����R)�����~兺t���n8�<��c��#��k�Rp_%�tr����+�EP���a�a>'R��QteHd���Ho�F��4ƥ�Q��DQ*��~U~'K&�3�T�Jٌ*K�#�@A��BJ6�ޱ���]�,:d��|���0®q��AR���vfɰ��Ǌ�����(�=[aX��z����@?�S�|�2Y�b��X�D`������!��,��S��1K��v�����y~��=p���X`x�:�1�����y�(��4^e7&��J��W$���O���ۂ�jy=�b�!�ۄ�n�0��4�5\�����(mH���*q:�1z�00��0]��ދ�r	1bp\�mΥ5J|�T��&�Z>��T�]��%o�'��:�����\h���	t�7m�����<Mf����vJ����4˭�HI#�M$/���iQx�^<}E�fe�3��Q�O9pmw�����,;����X|6B'�ot_�|�İ�UsQ�;^3��	����������]M�(�~4NGͱ��Af��A���������0�'XW+LsZ�f}=ss;v!5<�;!��K�-%�a񏪄���" (��cq�܁��s���n��6�� ����sXxp��2,��{�G:ȶ1iD���!%��!b�W2Sg�1�<�{=�k碋?|q�ݏg���c>-�~i��_L�p�#X ���j�odΎڒ,����>�L���=�����m�{;��7Bnp-D���f0G�� ')����
O3��Ƚ3�����V�{Ԋ�a��ܙ�n��p��v���%gϝ~�j!��gܟz��+�09�^�
��TdsE.�7���v"��C.�E�-���^�1)���"x3@l��
]ͫ�G��,�
��qr
���[c��mлRm��O�T
�~;z�M��k���+�`���ց�)��w���.��K9�"q��,�l��]"<,z�2T��O�E���oa�7	8�gy��wXe$�嶶Z��W��[|�����]2 @C��~$5w��@���-�-�t)�M�&� �!v����x�8����Q�H ��� 4����|����(�.��Ka�Zоx��O�b�ĵ��������Sjl��z�K�w�:gѿ�<�!�2��˦N��Ue�ǊFg��	��y�t.1��HOh��.(I��lbM���|U;*����$ ���L������M�F��������@���.p]�D7���z�L�f�HD ��V^YI�(�h"u���7�0�n1-7T#��[�Y����a�渜L:	�N�h�%����������7��u�NOj�E����Z�V����}0Fn��Y=!]ʶNj����nɡ��:3n��6�M��S�m�y��zg.��v�8�0���M�_3�|�I��pj�\XaK ���r�c������� XT+Xｏ��gx�z��W/�g}���<���eyIG�@�d�
Z�@����G5�pC��fAt�3��L�7�S�+1ɂ��&��nN���3=ll�g��-Q'��V��3��lFga38����R���ש�;��������D�9�z\4�<?*vH��һ�;�o��&�5�	9#q~��d��Q��V�G(��L���5�}�/� #o�d4f�Ϛ�wK���+��^���B.X����7���E:�:��G���UFs������59÷�����У!��}����Ѣ�P/2��)`>2��;�܀3C��a��O���h�Jֿۙ�H�h"A�2��z��j���
�e�QdA��!V�(D�������U7�^�~�T|���3���s1&���L��
�S$yx6� �5#?���4X׵5[X33ʿ���\0�o�+4����	M�|"�+��v�e�.��4�d��*h2��F��u�[�i�s�c�޸@�'�ޝ.X��.�SQ�J񼆛�¬�P��AP�ϝ���\<y�.	����{��n�c�t�$���z#��jt{�f�!��*�`�(l��U���>8����$7�NaU���J�~}�`�	��W�����'˩�-_�H��b�+��T19^�b������(M*Eo	r���T��R�����R��mW!w�S\�=3��[y����RM�"*���:��vO�����9>�j����u��`�����֏��4-$�f��dW�2'�^��l��
����E�k�}��Z��[/�y�j���\�:7��Na5�2]�Qxk�B����̘c��A�Ʉ��=��O���.Ԙ�����q]��D1y��<Cl��)'0NXա1���p74/=�8�H�ܘn<9??��{� ��sp�w/�FC��cb��vf����E� ���mX"��-L�u�4=e͝	���\`-J'"׷�_�2��ؑ����N̙qw����;�]ƩSXouT�[�סRjM��D?��cn������S��$]Sʻ�$E�2�EY�ʥpeo2���ʪ>� ��Ɛ�������+��1d������A��C��g��N^��x	�����\8��Xǔ/�W�Ņ�CJ����>�]�VA�P��'�����QStKr�S�����IM�$�(���K,�?������Y�p�f�+��dN�\�!���s�f�$�;v�-{n�R2�$�g�+JQ�|�i�1Vl���B�0IZon	."4�z��e�i���=.������氃H�?Ok�Cmg�|������ȹM"I��G��A&.}�.l(�[E�uG���HM�k�s�o���Zfߧ���O�o���DRr�8��X�Q}���o�h|��s��=����.�m�K/�Su���?}�%�Cנ�]��H��x���9˂�ɵQAi��H�c#�e��z
.P֕]U�9�F4���ѡ����U�jW��WwC0����jm,�\�f�W�^�~Il47k&TW`h�Q���:��^��;�w�^e�|U��\�fe<X�O�>��W��FQ�w��rh�F���EA��@`|a��W�I+�����?%�����+�Ð�|2ne���+Y��߷RP\N�ݠ�X�ސF5���I���o�3�����4��-g��ottZ�[J�mѼL��}s��8�3�p�Êc�j*Q?S� �!��#���6����� �H�턤Z4���uRO�f�G`o��-N��������5��x���,�R�<�����vC���0�7\lZ��G���F�iq���
�t+`O�Ñ�_�q�<��#1203y�q*�4�7>L�mF>�$0�:~�,d�/���P��s�AM�?��P󖺶CP��K�N]P�i�kBbO�o�`�h"P2G`�Bi�ى�9"_�X�@H!�<��6򦾴_�[Y�s��	,3�ţ�=�qM�L�T3�)ZYwlW�[G�J`�'v� ���=��cz%ԅ�|\����p*�cf7F�,�T}յW~���i98ڊ@�q���msM��U��_��)�L��K>UȨ���t����5V'0ZΚ����
^��/�B�a R�/W�a-;�����y`Q/}���Ef��e��VԐ'':�M� N�����4w��	p#�.�H�˸�E����>�9��\�|}�_.hP�V�� a�Nm�ᖡ.\�G?��}�L�نRWҼtP�D�@��_�Z&#��yq��ч;��	��<Ѕ4Hk��<í�5Jo�~*�_���2=�){\Ԁ�R�x8�[�N��'���"_0U5eae���m����G��-��k������T�k�-�T悴���C��g����Rp"^�بϷ������$��N��v��؋P���3I�%z�=r�vsw8����]#�ۦ�]"UFL��<�� ��/�R;�Y�@(4H�
�h�̍W�	����
R7������It�:�VR��ʾ6�d�����b�˺�n�=7n�d�i��!R/$w�v'7kL2���g�Z��K:��q�Ws�2�������'�	~�V��	���v����-!��a�������*P�>?��\b$5�3��eS��~4ǁ�6�a<"��'�#�f�E�ϑ~����Q�8����·A#Otow�+��H��+�7�݆�߉xL/�gf�
c��H�Z �sQ(V��j'H��-�CX�y&
;;z�(�(�J�����>V5��M۔�ӳ��A}m�լ��!��%am1}���]�8��:���S@�PD�|����	�Kn���dHe��3�q��!A���7�(�cg)��$�M�tT���X:�����qq]Q���i�/^s�D⒏���bu��uN�+��3��0�z��dsM8��Dz�;�����#�efl��E���o����O�ʈ��~:9�곇��)�*i%�pY���%��PѺN��r�|V����$�2�`Q��O��F�������1��x�2�K��A�~0{I�(��"�!�G*����KEE�[��o�i��Y�ϊ�8�`�W���A��Ewu~�ʗ��?����X�XL�9�BYjF� �C�d�J��܈��X.�1�8;�y�<m�y�էޜ�5�$�nX�'d�D/�S^�[���2�R�W-����f󔡋�����xZ���oGj*��]!RM2T&!=a	���h�ǯe��=Y<Q)�_��%v�ᆶS����a�_��Bc�ӀM?��j��[Cn}�	v��X]���n�U��K��a�|���?Y�o��)|Ӛ?�H��5�_��jW0:��y��7��Kw{�j�޽+��>����:�/�<��Qt�]�)	�����(����p��Ek�I�:I�]��$�Ug��|�2�uj
�m����J���Z��bBh�j�q5��6�:������+��/�����G!�o�^J[sy����/0��QL�ul#b�����GHZ���f�Y("���5�6RM��7��J��0=�6�VR���F��{O��*��@��j�<��|��3-�̓d�K�Z��է �?SY$�.}�)�a`������$�k���ɚ�.صG��d��
����2��s��I����+�>B(X)~2:M|<["��C*�H(pL��s�:���[�`0�����!�����+�}����i��Z��z��5�g���g�1tN���4��x���5A��$=�!��	���e�q���Ħ�0.��"@���:�eb�{Ǒ��JL�ʻ:��5O������MNO��V,QD�$�ڹ�}=��|�ۊL�<�(�E�����{��ي���2�h���M�-:�U
c�-��#n�x���T�C�'UY�T����9m����חH�����Iڡp�u�B=V&RK^�������FYC�ZHd}Wi!�d�{�OܐA)�V�2͖�Rh%:~�_��=��C�_�9��M��M��>��[q�lE�0-�::�3��%o�vN�q:n�=��Y��&"��F���6d��f�%;a���Zi�gs�ʈx�֔�4r�����eh��L
��Z���Ѻ
bm�}c��f����+�Ŵ���2H�B>����'���T��=�p|�����%���IŨ�"Q	��.ޮZ]��[��}���i��كKd!�y�,j�?Y�0��n��y�	�{�&�wx�l������{	��}al�r��n��G	�&[��|M)}�>J'�~�����$S���ݏC<Bgh����',��:�:����x����ɺ��"^3u�]s���=g��oo	aO��}�"��K�+ټ��¸π��,�hѴ��%�ڠ+�7�����RP� ~�+�-��2m�9)�c ١�����x��U �#mϟ��8�d��&�,�ϓ��^�c���/q �Z�@� q�x=�a:�v�?�<��Y���,#��G���)"�!i����L���b�`d�6'�C�3d.�U��m�0mU�a�FAu�����C��)��rz��Q�	�������$Vc��|�ޘ�o[T;�)����d��jcG�[�g�ҍ�R�˄�����.��Y1v(k�����4Ppcn��U��X#�º\Kٓ��)`V$�\ķnR(��o89T`Y@a�Xs��O^��C�Q6 �*V���f�~��3Q)���z�%�/TMS"3a�G�$����I��a.�sq$Li�0�¯�S���I%��.���|��P0z�����M8��b���<�9�g����ԝ�ԥV��i5�ly�����H1�AJ����X����Q�����>p4�:OKd��W�� ��H$��?�n�|ڹ���n�N��3_��>th�����@7Y�����Q����d�}T֐
Jr�5��&��&����bP�w�T퐗8����q�M�Q��!��C��e����a�0'�*� ��|��x����Soz�HT:H�fg��t<;}�NϕL�ҵ�[ҔYkk��c��Z'��bЛ�/JDUv�|�e�n�2���Et'���������/�)�ӼE�v�5�%�y3+�8�-��$�k��t���NF h�[Gte@�αH�AU�wh�q�H���p�M4Ō,�e��<GJ�x_dQ�0�Hf��Ij�BL��U܈�޸Rv�<�ǋ��ơ��g�`[��gU�t$���90����x��ĺ���\�,;�v�-qE��ݷy!�eG��� u²G7a�1f�yy�n�=#r�C˙�b]@jg]�~_.c�y�YY�"C�u�+�~ß�Jm��L^{��}�ox?W�Ǡ2��Q���N�Q�;���e���i8}�v��g�U���c�v��ğ�2"R�/���S8	x3]��EJ|n��N(!Q� $(�ҫ.�AH�T��fl0��%��#,�z�!F�@9yL�w������5{,Dz��!�i%7�b����r���̓�3�˃�!�b_�ox����[�SW�+����1.X�2fe:��L:ȇ^�i��X��ؙԸ�u�y?��I4m!������}����k��| ���\GJ��/�"�NY_�	���RMD!/eO�a�v%�{�\nq�p|ͤ�,E��,@n�N�9�.j߭|	���z�P>�X;��M��C?b���`%����W_a�W���ST�]�-+��y�d�v�7v�����f��l;��a�W�N�g���u�BjJY6�S(�V���9�l[��s��Β��=/ۏ��Y�EVw��R6'E�cɢ��e��m_�ϣ���`����2�$�����>V��~
�N��������Y�`|B���B��C'�ˠ�'������*J���U���h�'�9�}띩�'z>%4-����j;��;Ef�Z�������Z�
6�}s���<l����]���EQ .���g>�/���M"ǂv�r�'"Mj₍�b�Ne�&W�	;�ȇ��=�aŃ���8/F\��I��8��1|�=M�>:��0.�[G3K�8$�x�jdsã��#jن�uUI��E!���Q"z�q$r
E_���_#h�g���S$�@]�-���OɠJ��!R0�-�le�#9���~*��&��`��lG��'|���G@�h��):�[E/e��_n��mиP�Y���M7��d�=�.;@�=P(�w鸠GCeb�f.P��)�$�S���ڈ�m����P�#!��ˈ��k�G(Cd��{���)ˈ�9�n7���V���W'L�N�w7�����3�O�òm�g�<�k&*��$#�A7�eM��M&iZ&L>���Ux�e��á�;(�M�̓�ⳝ1c�� }����X\����#�K�˶�pe�g#i-�-��}�q�'�v�f�0��W�Љ"���������������GG��؋�ZCSR�ׂ����R5">栖���Ӹ��.M,������K��+=��ߵ����p7�G���Wt�U�b�'فZ�4j�Jόt��T�=zU���ꯄ�ؽxv�{[Տ����{��(�b����% �� K�憀v������.�Fnn��m�8D�;r�f51%-��
T�_2�:�p�b�u�B(����g�s�ܛ�5p�kŢ�ٕ�P������T~ѓhu�%�n_�8@Y���=��[��:�X[̹Lw=0Z������Q�"�y�����z�:�ye��:��Ե�'���PkOHW>��j|�ݪ��\�=�5� ԍ���0K0 ��Y(h$N�ſE�.J����g2��ajh�<-��| Y�bᓞ̬@�y��
���мc����Bt�C6D�=�s�)p
g0��,c�#��?��lz�
e��O+L����n�� ^�V���(u
����x�3Ť��S���僎]>A�^Qaۿ�����u��!��^	ANd ���ySf�kL�S9����r;����GA׵��u RZ��4ǲ��衻���Q�_�5rl�*��f�zAᙤQZpk�� tv���o�(�:_f��v�{���)�
���;,�����_�,1o7��������:3��gs�km�LW��c[�aB�٥���������@��_�4j���bD�Xy`)5%��}z.�wdwj�������e�4��Q\�5ܚPe��̵�o�8�?;j�Gt��<=i^g�������j�+��(C;]`]���>Q�*� �A̟r���坓3qg7����]߭��[�<��z��� ��7�W�:Y��j}ݎrce��k�h���06��@���0�>%dqm�RM�]�[{AKt��n?���ԗU��?C;�M���}9�J���xk�������[p�@`8����-����J���R���ng�j��?h�7���7���Zy�4��1+ȗ�����-=\,����j�8���dh���� ���H�ً/���_�\ie�M�N�v�ꚝ��F�+Q��<�]fZ\��8��Ab݄��s��@���A]�z̘,�*lO���ŗJ�[g�yW\-���[�� ̆�} ����B��Z�qe0�g ���	6E/��ǝQ;dx�5�k�Eo�|��kL�˥�l�9�!+��|;��D�.�V�̃d��bN'�M�}f����&�\���݃�ԯy��?���6]q�C��AR�̋�<�F�b�p��>R\�X�!�<?N�W7_�����T�����{���>O;�9Հ�>n����K�
R��7!�y�7�O��+�����r�R��Q�VY��=�І�e֖ش�wt 3��@�d����"�o�y-�/�q`��]\�<{���1��ʥO�����:�w
�`L�}�꒫�1�<�3��E���]x��O/�i$�S����ls��vG;i.V�Ĝ�Ƌ++&h~��E�G��U�>w��̳	�k�6ک{�A��7ɉ�}�u�;��%�Ӯ���t���,y�d�%��A1?u7jo��J�_���C�g����a�0��T�'��@���#����&J�S�m-�
a��c�Г����.��lh0{��"�v�F���ĺ�(�d�|`^��k�Z�.��^A��cW����;��|��}] O��a���RGQ��3������5ob�sͲk4j���عk�.G���lU[���[1��n��_;��U��0D��a׉���SL�1B�ODt6t��g�LN�^-(p��z�a���m���q�^{�b�])o;��w tk���zP�~�Z��,��3�@S��B�y���5��a���A� ��|9*�z:u�Y�䒢�|92M}�nE���r�>�5�c��T?A��Q�o�����,X��~绅��c~� �G�]q�7N��^u�&>�Y����?�u�ER��4���fۅBl�B8��`��{(�쥾�����pF�+UT�m�xE"��שׂ���0�=FJZ5bƹ`Z�[.���yE��Z���?K_b�� ���'I�%���F�6wH�>M�}����o#_k�	TC� .|Ҕ��wO,,��
�I�l^9��o�Բ��!�t�ȗ
��E��.s�P��?�7�I�H�+���lh�?k�g��0�KQd_�i;$r�ˀ�/X��^L�!O�?h2Z�0'5:���v�O<���y�"�U�e�1���@L�~l���ߟz$=أzc32Q�2مvJX�O�~,��{������CW������e����/����[�z�LI�ΤP1~Z��t��-e�,���%����}�Ҽs��͋���&3�0̹��BX�G(�
�+��z�n}���^��坵�nʼ����M�m���.&Lp-�#"%C�WWT�5�JZ�ŭԨ�%��f����^^R7ͅX�"m�]�o�C���c ։$�L�;�rK�a\��i��ζ<��w��)�Gښ��Gb-Q�G�E���aT,��i��1'<�g ������w#�ղÊ���?���wo/��;O�g�g���`��	br`)u�[�.ƌ�4-�W��˾�5��Ɛ�IQ�P^M�t�D�����a�r��;_�Z�s> ���\� �w�U|�������~bP����m�떥	��+�2��7��ǈ�}ǚ˞����F2��r���E(f�(]-P�&*�x�iuX��/}��:Ćg�f{���K�Z�yJ�q�����4��}��L��E�I�w��֣c��+�̝+�r���>T��+��,��<�n��P�"�eu-���[���)�,Iyn��@b���a-����l8��u�3�Z�:���Юذa�o�
�052�}��o_��V�沁Vՠ�}4�sU�+wVZ�?��ȝ�[�!�E��$R¾A�3��kJe�j�ջ����2��V�y3 �s���"/U��,�D. �ꐓi��(��C�8J(3\�7����"}����cF�H|��<���`�#�|.��g7��}��T��<z��e˦��ł��5����f<ø��ܖ����>(�-	!�_+W���	�Ɨ9f�P(Fbau�ݍ4�#P����~1���/��Rn���֣�a��,	(^�!P*ucN��iJ����[�V��W��~�IzBz1��!�Ƙ��*R�N��(K��t��k��S�+gK��V�k�KF+
0�N3�r�/��"d����r�}�W-�)x��Q���U��#[��|k��^iJ�<j6��{�j�bRp#�7#^#ǩN�� L6l��J3�*��w�����=19��R�|�S]���!>��؝����\_�]�_�(w���KG���Sr�a�|D���0��ݪ�@'T�a��5���������n���G�-��i��dj���[���5w���֩�0�d�Ĵ ��,������������ʱ	p%m�K�;�!1���ݬB�c���h�%����d�?�&��*V��`�h����D`���,]�g:F�':���n�VԊ
gl��D:���=)�f�%n�Z �ur����<�[�ԧd�->����l��wf��N���e$bf�2:�A�{�I�,�u}��%�'��ƿ�22�9}j?���\��hU:��ɗ��1R�g`|��vS�c��0w��6+���pRB�����Έ�ܔJ�T�Y��{dK^����-2|��fBZ�9���5���>��� �:�8��g��X�ߤ�T���xzu� ;����d��^���|�x����6�I6��o��"	�|٢h���c�\l�ru&cԨ����;;}������"6����5����£��$i#�Gǿ0����U�wO˖�H.�\��1d��#\?k�Y�w�(-(Wղ;@swL����۰{u4����6� R�:ΦkƓ��g����趬�Щ�7�����[*��~����H�	l(fY��R�i�O���h��=���o���[���-Tu�J`
)�������$�~؋����f���Ł��¶@����W�	�[j�f!т�r�8�Q�*s���
��o��\�������
��h�_��� ҹ�D�d򛢜T���d�� �>����A{�u%ˌx�|��������m�lN��>�͎;�8Eœ����'w
$��x�?e
A�وxҒA5�
�����_R���k��d��⍼�����MX��'qk-�U�4|<��2C�.�ӫ
t�-m��
�^%ӝ��oߢ�rh؟x��M���bPc,?֕�S-xg�w�Gg/� �s��[��VG��)[�~H�!�g���@mz�z�{ ��!q�m/!��t,��/���v��4�NG5��}�9;?fxa�_�]
����z���u�U����?���8I�����C���QM��r��ʾb��q����sCPE*A�AQ���}12�}oi	��]&�L�`,��$H+#eʠ~;X���g'�1����Ū0����OV�?noeD��o�%.�P�J�l���)#H] Ej|����VQ���={�����게��uĳ῕;��B`��~�)��׭�ļ���D�!��=���N_�e�[�!�[����)�º�]�p�\�Ml,�{-��1N~/KN���Vw+�+���.-.��M2�d�_Fc���WL�Ľ�g�n�:R�B���}�I-��:ls֔�Km��G�۳���U���4}Z��E`Y��vK���x�+���w���:����H�n"�P�&��*�����%��୯��vv䬥b�.<�}�`�������7ZL�ﻘ�W�_�x���Ώ>pB��@۪��ۖ��}�	�C��URT�����(���:����ֵ���(HQA�ۗ?BK"J�q�|��i>i�`�M�s�����:���UAa�^�ё�,T?��#[���E4~1�����"o��U���0k� �hPv>N��ᰌJ]�~m�5MGX�)sM��<�W�"� 7��jϡ�"����)\q���ڿ��g��Hc�cw?"s�os��ϡ�Ţ��sB+Cn���J�
��
�d���I���R������q�&�9A��r��!k��OT��3���l��A)���H�g������O�0��u h��g	��]Z�C	�R�n���o`�ڂ$?���v���I�'�2������_��ml0��%�_f�/��S�u�=��2��
��e�Kpz�v�XgX\
"�@�2H���^Ý[�
��&(>��n��!�H=�є��Udн�⸟���-���AT�[���=V����&�.�щ~c����P���,��?�Y Cq�/KQ������J����G��oOp�{�?I��4�pET�~�,.ݍDt�ߘ�6�S�>s��L *���0�RL#�S0Jz�h�,qQr�����}0z����*z�8��y�l�}��%3D���
;��$c�^�C�LIu���Y��!� �-)�jJ�0;���F�b�C�:�T(!crs�N�
G��� !f��L�2X�uK�5�;Q��.J����.�P�S�,ŜK�f�fm�gX^��<r(8�{ha�[��Rx��	��.ټ��WT���&i�;�=n�>�y��`�3�uyQ��^����>���D��)>��@N����P6�W�*����/�/k�1���ը�^u�5������R��������0��"�^�!:>g��S��i�Ő;�"+ c�0�����-�0�� �4١� �x����IN��g�ఞ+�F�F`�Lb0�WwM���$H�~���� ?���EH+�ʆ4R�P�Y�XA �
�G���/T���Yq�O5�B����XxT��m��jwt�%9M��׌tu�<z:�F �dL�փ/0�|f2���v$L[%G"��#����=�9���G���.vRV[�Fx0�hu,r���z���TG�wu�}Tn+�����+��P�iw�TbDҗ�3r��u�PL�u<�>��#�#s��E�ȗ���fH�	WX?��e+��ϖ���V�3��T�f[��iP�yI�T��8�����)�M�����|�r&����4��>����[x��cmD�X���mR�:�&���U.��gR6�����HCB����Jz�I��e5u��K�S����E�qpn�8NPAo�Kk�	��d�μD��|a�4�"��d# ���\ ��x)���@h��t��x��Gp����C����эB��/�� O[ں�4# ���b�am��1��� �>�eu���!����l�P�WSM�e�K�5�����3ln3��A�~Zb�R���h�(�I�{���E�l��\[���}JPsɫT�q��L#�X���)(5���y�vӃ£,G0���l���V�B+:t��4͐�y��,k���h&qwm�ף��8d���sL�Ή:W�Q��L6��,���٤e��L]���Ƃ)�;漴Zp�]�F �B���n��y8���Em�c�h�@�}�듨_�-|+�t�'�����P���b-�}�[Q����YG�̦�B����f�J��^���';\��݌4�f�=�&���ESy�}���4M�B��*a���y5�ͳ����
�������m���R��v�#,�������F����̟�9��HH�ƽ��� ]D3�"��=���p����e�H�N�/�dy	-'��L�Ψ���t����#qv���y�á3�؆�gV�yۘ���.��D3��uj�q��8��!H^G��C�ӀQ�{6���޶
���g{��c��E�MQ0�Z��f0ķ���u�̟�wȭ�N��e�6dH�ʊZ�,��I�7g�M�<�:㻩�B��PB������C&^;֬��eQ��4V7�0Ugƺ����q�-
(��z1���u�ָ��yf�|A���ښ	U�7��<���#�9�l�_7I�P��f��a��3���6�~������?U,����b>���������2�m�N��U���U{�s�}8I���ZP�^�`�����n���/D<r+����,�b��/6"%{�� ?�U��z�	� pу`� �o[�=X+%eP~�W�sk�L�z�[��(`ߒ���b
X�վ��I�-�?l|�| �m��G�y�t�`D�)�횗���]��Y��\� ��f�@Y�@��ޮ0�S�h1=�"Ha� ��D%_��	V3��(7P�[��l�r�]A�(@c"�W��������PSܘ>n�i�r�4ތU�`�q�(35����m��i=wnhI�d>����g_���|��6�۴��$�<�g�w1����œ�Ux����i��8�}"礁^�tJ�Ƶ�T�p
Y�l%�mp,�QY���p���"I�����+�CٍE����S��aL�� �]2T��/*9��������p�25kO)���Vg�k��\��~�J:P�A$�?�U�����J����P�����dk�Hz(�cs�OdŔ��bn�*� ���j�t�',� �ڂ�c���|kO�a�!JB>Kl��h<b�O�z&Φ=U�>y&P�Cv'��6/�O�/	w)$U�MDaF�~�1`QI��P�?'jb�#9��(��[���
�[���U���/[�l��ԩm�1L�n, nҰ�ɿS�v0��U�����^�(��*�.��*�AC��Z�!8��:VC��ß��o����
��	sR?��Rk #E�l;�D7�ҕS�N%\�*S��a\���]d�^;}x��<b�ZG�:6}�^��m-��ۦ7,A�I�3W�����&yXL6�;4�I�x�ەX4���������܍$�l�KV+�%�/��hps�R0�&[���#�hp�����x,ﺷOh%����u�-����#!�FE���S��]RUp��\w 	
N(��O�F�+��z�DM^Њ�.���À���'{,�)d,�iy�Ǝ�*�s�}j�E�S�|�����W�&�<U,9��[H(Z�=j�J��^� J��b�]n��*_k����ٞ�fvK�hY�kBf��-�̺1�f@����C�ܳ���:��, �|��KŗL�L�|W��"�j�_{����f�B1^�x�F�ȼ��&<�~k�p�zy�e��s��x:�[l<��Di�3���A��$�f�$|��&�x;M�X�O�^D�a�cr��(�c2q��C|��e�=}�ۿ���ușf�1C��BZ#�oMA��Tj�)�����ɮ�|�ڋ
j�Z���|GМ V�xO�.�=��w���9J�֏�n.�����W��X��WEPܐbN��%E:���)�^�'��zM}{qt���Y���S�t���XA��O�%��J���г`؂4�fR�ߨ��P��ɿ��8����y�#�2l�SLy֭���p6:1p�7q$i�O���BK�=�p-���
&X��i��W���j`ޮ���A�d=.�C��0bjn�]�߾�Q�*�UZEt��Q�و�Z�Sȓ%;#=1AI�d�O�Xr@6)5y��
�K�}�"][@oiC�]t)��]N}��6��3�n&A�2�W��$CC��6*Y%xF�$"l���CU�g�@gNֹ�?47�1��ڕ���	�lŗt�r�*�ޚ�R��w�2'�Qw�ϱ�F��v��G�ɀΥ:�M��8�?*׻�?�tE����6�S�9�K`V���;�"��_H,�'P�'���vfKj��LW^i���C3]l��A��B��R������_hd7�W���=o��!�� �dd~�7�ż���<:�79��9�.����.����0����Xa�`Ga�R��6MJ�2�˺���t$�`��3FR읡��s���hi�Gfa���p�k$y�!ѡ0��,]w��޹"�p#�ۊ8��d��.�[��KE3��l���4F��6�Q���J��P��,ѕ9l(膟��c� �Q��Se�s�U^<�u�,'Xd��]�\ 1m}�W���������r{/����N�X�n�ڥ�S�/"������h����jd�
Շ5���j�<ی���8��-�X�f���r%
�ݧ�? � (	�,���c��!v�w�i3lg�tmgcK�^��4�zZ,�&����RZ��qn�� ��B�r8�w����
q����GJ�1:��Cw �y�8�{m�w��P⤝�h�)m�wJ�l���E�����~���	i������zQy�q03ї�2N��&�2�zt!X��AU�D%����ҔLƌ�=�Y-Mx��/�y`�����`�� z$�j�E���� ��sY�@Z����X%GBʕh��m�LY`���P�ӡ� S;��.��p3b)蝬����E��|�T�7q��5���(F��l@������ո��O�-޶]��s Kg��g�7�J�XD�r���-M&�P��F�~����17�f��Ǉ�����?.�v��Lt�<J?9A����ೊ���PtO-�ld���צ�����P��oo ��F��j�G�KS1m>�@5"�΁�*y���[��#����c�݇�}Z!|�a���2����a/э^�,x�A���3��vH'����-��z��Lܓ�}d��U�4��߯��Ӡ�@E��2oU��0S�!�Ʀ�ch��3�m��K��I�
H�*��gd��}/�Ո,�����oM	���:i-X�<-�*�S+:c��xJ�b�@��MO�j17�W��y�m3��$�Q �{�l�svZ���og.tL �0�~X�Kh�8g>fQ|�X�$�XG��
Ԋ~��i�����h���NV0n=A��6E�ݧ}�<,��E�scf������;J�P�f�{�f�=F�]ɇgop��D��C���RlMb�5�WW�U	�{��x#����W�%���nO< �Q�d���p���c�\R$�������x �f67� X�v��4y6�^����p\�=5�; ��N�Fv$�:>K���=����pM��B0k�y�˚�L7��N�VL�@��H��%re�hn�I��c8�u=��)��cx=G]�����s�T2
�<����p�ʢ���1�zD�Z,X�7p\X�;�1V��y����z��f1�3XG��_���WV�.~�7�2����������@&;��}$FL����ª��T5h"�D��pq���b^��c+�\��o���_%7bu�6���q!k��N�W�A����k�QzЏ�=�5`хt�G=��RQ=X�A J��|o���� ��+�����＆@�R�6?i<zѯUO�_&p\;�߅\�B@��s���t (����L}𩳟�͎��2g��Uݏ�����ȍ��}�:K{�����*4Ը*����{�ʠ+�f�M]i.�A�z�.�h9T�w�1_	pWw�զc�~��ެ�N�3�����E'����f6�p�E�������>"�t���d�OH����(��yQp9���*H?�ah������0������S#��<]�x.P�VC��0���i�����W&u�NƝ�`�\����W�J�W�]'"�Y�N8�p/���I��ǐ����+;��`�ӯ;[�	x����f�27%}��:v�UoQ�Ն3�`���6&z��b�G��ɖ��t%��>�#D�Q�\b�I�	��C2}"۝�xOBB����g�Ph��.����Q�A�%<N���}��G�>�<s�'܏J:�t�u,#�J�ߦY�,߶K��'vD^]F���# 8-�?�3HZtŐ|ѵ�tKq�X�����B���h/��T����q��~����@�]2wX��3B��;���0�%tL�ѵ�ʦ�;�dҍg��~囨b��%��"���"0
�f%�v�&	gJ�q��������P����!P�����=����݋��U��c0���£_;A��J���N�6����K9����oѾ�)C� �H�Lmv�<U8����yr�2��I�+D7\��d8jmL���gW\zx�� �Y)z�6>�|A/|��B��I�SX1�q��϶_�"�p��8�����Z�Q4e��5L�G}�(7�Q���ɞ�vvi�-�`�����{�^|تS�/�mg)�¿�8h�����A���^F�;�p��W�O<��5Y�	�=��F����+�'��g Kbڥ��e����XM���K��}�q=������le���li]g���~�{?�LB.����h�Pe,�Yi�k~�qL�b��T�h���W�g���L����J������nu*�7�����w
\xK�.45A/#F����ܩ�PD����7�x�X3����-��[4h_�H����4*el,\�/1����n9��;6��n�)�8�2���H5"�Zo��N�y�t!���\Ȱz�ʱP�OŬ��\��)�/�9���6̈�۷�h���"�/�G���^*��=�~;*Ĩ˚:�Ģ�j��^"}:<9���@- ��]�l!�g��Ta�*����Ȝ�e@���׸���J��5�ʽ6cD�f����
\�� ��J�PɊ�}
�%��P-��9C+/
ޙL�=�!z�ひ*>�<��Ȧ��)�p��lI�"\�~E��cH�J3� w���`PZ	5d�4$�R�Oōs5{��R�\u�E�NJ�%�& �;�;��fz%�H�"�d��EQ(Θ�Wzu��V��M�D$,#���1M����+ea�N6�v��ْ�xYV�I�9���L-�tK�J�_�]�w6��'�ﳧ�%��Q5��Kk����Y�	x?�����45dGղ�t��T�G�%)���(@WH$c [��G��"R����,c�$IP\U��,�7<�tr)�4�rV�i���ȝ� B�-nc��J������V�ܽmo�&�*Hs8r�3E�0���O�eD����$T���H�$�����~r*kz�p5]��`��l�>���Hx���J�C�n��׮������i� �����,�"m��7G�9v�#Z���B�GCȊ�lEm��!��4@�aKS�/�Z^���I/M{�;G�s{U��7	UT���������3d�-��,J�Y�Ku;1�2�-�Ϡ��2Qx�X@��[�1�Ao�ٖ:�$%�P]7�d�|a��4��Io�팫^qd��+�k������*�G**�n��=�JbFԸ�So��$ѓ���;Y�g��7�Gd�\�O�-Ώy���ߞM����,m�/kY}�LP�a	��]��T�t�	��r4�n��G�&L��9�խ�>}���-A{?�;��DV�>�]�N%�ow�`}G7�'|��Ͽ��b�\���8�k��9�����/%�|q^����tH����	Pp9�-i1$���F�zV��c���	�}u�B�lM,����2^�Z)����Ж�x��J�Nj#L"�^�Я� ���H7�r����Ƣ<��X�v�
��G)���_�ɗd8b�Swa�(s������QuƢ��ù��8�2�̉q��(`lY]!�G��-�݇~z��x�t�Ⱦ����y=^D�#΄ڷY1�r[^Z�}AFg�Ԟ�?��j�5�?K���U�{���s�-��Rm@���c��c�u� ���Vy�N
�
��eC�b� �lJ�$
z�J��Z�>ϯ�g��y��\��8;f��Y��}kP�3Rm�%: r�6sBp,��lɣ�=7��cG!�������BѮ14�zX@�QڷM�
՗��֘$?����j�Um� 4fT��P��ī�`,�ĝ.�:'X��ԕ�ny�m�a�` �%$d4[l�������k�ki;�S�m6��狏��8��)��s�j?��m�԰��Œ�ތl�VJ�^��幸��n;*��Jʬ�����{ї�L򓌋g@U�?G�e�"�oƢ�},��WTW����}4ykt�|0 �o H��Ð���c�`!MW%^�dG��_���y<S,��[�B�����'����T�Pw�}є�������Ǫ2R�|ҾM������P#2ux�rd+�U�IZ܏WW-G�a{.���B.�p�u&,�UJ�ȗ��0�2�g�
&��%�W�GP����6Xz~|�����_�ٔ�:�|�7��-������|E�;�jԍC7�$!ڟ�7:
Z̎@�nء�p�}�'�׭ϧ&+��H��g�L��L�	���)���)FG��	��f"$JjϐK��������:Jg�������ng~F�щ��>�*Q�p�t�Y��6���c�����U7#�uI��)�dg�B�p�'��%��T��uE8_qw,n@p�$������Ah�!�_p�|�0`�s�y�WU�2�=Ba%��q,v��+����k��堶Qâ�i�Q*|0�t�Q�n|��]�@��A[�O������F�B�%�ԛ�Ź�B��ɽq���[0�׏�2]C��4kC�P�}���G*Z+W�Y�*?S��Q�I �@@=���>)0�=��ƦfF�L�2�3{)�D7��z�;�q�q�,(0��xyu�_@m�JȺ¦<Fș��,X�Xt��F��ny��q���{t���F�=�5�&K��Qn�����ꡠ<��_"��*#C����H��ITQ<'�Fǩ��̭��a��D�x�˄��&a1#�?���+	�w���h���T���[h ݋:�2�M�B���_���t֤�L�H���jl��g=�,R"��ў���FX�7~ٻl1$�#g�I!j�K�����̪�l��Z��%x�⤮���� CL)�� ?�}Lj��zTאl�;�m]���tu'@L\~mAn�R�tvn�x��m��腹��?�i�P���M��7�bC��X�=�������jϠ,�@n����U�_}�!$�n_�\��ި�/��ٯ��VLg�J1-� �t�Fc�u��/Z���/;�tU�V: ��V>DI,0�T&_�Xx��l��Z��� �ۉd�����Q`ڥ��/���`�V��apר�Pۿ6vYl���G���0�����V�6t�h�!�tX�msE��e��}*Q����o��~���H	P��$ݎ�y�Qpp�ҼuM�'C
�,~���J��>��6ۺt��ˣm�x��3=��a��_��b��ݫ�kq�B34�EayD���l�;#k�;E*n��݀�ց�%�1��?�7F��o7��gq�[&b�`��Uh�g��E����Ycu|B/�ۗ~��)�A�}�h���94E�4wƏ�wO���Il+B�p��&B��M2�+���)Z��vp���� �Z�"��-	3�����rMg�,���Č�u���1�r��Wm+TO�M�w��/���aj�@�A&붎��)E�%}G*�{Z/�ũ3C��}MW�$���$BL��ThTH�oK��GRo��f>"�{�c��F�o�w�����N���_e�۾���@�O�Nyr��I	[��wjU�nq��
�Y��ٖi.?���(U �Vq�� Mc��`�e��H�-�ۢ�����|�g��=_�%LQ��C&�W�w�pX��x\z)<�a�&��%�.0�Y��fƁ_�δ��|aҟ;��ifU!G)_�6�Qu2��>�0~I%{Iu����g�5o��k헰��VD���-#x��׻R47�u��˃�$�Ŋ�YW��4"I��R��ɥ�p_�����]Q:�xr�O�%U�P�)cV��/��l�nǿ�� "ž �Ewhm�aUc�tuZ�AY^�pK��@��ݡP�i�'{Pї#��@�I����\};�_��%?ӭ]+j��yTPz�	4g�_�D�H��a��^z�
��-sC�P���Z�F���2]��NJ�����u�}��N�A�:�Յ�NaY�wVͿ�e�N4}����p��j^��K�%�we�ˮ�v~K��'o=&�/LJ�@��M�5�2J|Y�lg�p�a����gǴJU�G���m�N�I��9�^���U�KkO�WS[����yu]�z����^��+��|��2����{�@��0�9��)K�5���hԭ�����D�dSV��a|�Z���j+4�Z؜�%�u����^ͫ��/�;h��ց�ks�l�k��^��2���������+�b�!������D�?��N�3�o��n�a�赑�/��&�@��l�$��+��b^@T��~t�sܰ�0��XVun�W���3Y�ſ���\��DU>��yPG�C�0�z��dN�j�e��1���!s��ٻz\H�` D�iVo*���&��F�:e��� �s�!�˰���)Ӹ��(R�\��Vf�pʃ���;���^j=���Y:`�,�8R�5&j���+r���j/I=D��<4����<iB-7��^�`��c_� x9����)[���B]-�@�&�k'�W�MR9$�Wo��I6e;��f�^�%=�{=1��J^y.Ҿd(�0�m�g�E���!p>hmBV�]&A�>�d��&�L� �Cov�n��+���G����c��ۭ��̚�^�$l�}ջ�)�,k+���A�,��3.d���I��������-�|]3���)�~)ޙ �r���j��j�E���%�&09���Êq�cM�*rx��s��V7ef�����X�!f�gkEBX�inj��,����d��a6�q���'	��q���_��%��6��gZI��Oi��͖0���B��(��VRI�%���@yL^���ġVh�x{~�0NP%��_ܢd%�� g����h�C�d��\7SH����3l���"��*�n��l�GP��{�`��������;V&5����?;�y%E��l��Tң<�����A��px��h�Q=�����
���]�~�.�2)�tǗP��9�B��X�C�^y�[�Jz��/ּ����# ��e�����<�����_��[g8�8{���
��H���&	��Y@%a�4	?�!6}�a��?c�E���5�Yٶ�0P5,�I@���8D$�6)f[�vx�;*�c�r^G�W���g�����F�����{@`�cF�+��T�Z z� $��:`�#`��7PY�Da�ni)f4���L��@����xǖ�;(,��g!Q ,�Y�}�Zr���ړ��b��p4ܽ��[�Dӕ��������|�(�7a=]��A��j�tN����j6��NN.E�(�h��i<�efk���4M`ʶ�{9�%�k}�Ұb(�	��"��Ҵ�͈y_�{I�aYq!�?*��,���k�}�\A����A:�4���G�Ǚ���\^O��>�s����,�>�ј�o�	������}dF[�<�LZ�R�9�N���!}pp����1����.���[�w�l@��g5�?t�΀���%4��ו[*Eo/�J�DG_��|�s��b��5`%�2�~�)�3t��tԙ"�1D�T#Nl��@�Ã>-O�vr��&Ƶ��K�!m��(�C�ܴ1�p:,҂y[��Px/�줗p5����s�%�E�aOUj���������#ŵs6��G��R���'N�	��u.���׷h3�b�O�@�hwB� �������h��}�l��"����F���8�<"���)�ܳy��9,z�S&$U1?"ݛ�)��CqF�o��
	m����P
a ����m�U�{����<���֭��(G�:Xr��;�L�iF�͏fm�tf��n�^#
�'��]��	њ;��R�a��(d��r3Z'~I��*M��ԙ��z�{�Y��h��s�[O��Q4�H�%a��o��3��V�u^���Qh�����zT����Z�~yr闡zP �)T�ӺO��o��	���;�_�\n鉣��#�xldE[y>�l?�M�t.��[�+n ���m\l�i��+:^�j�|������~*��%��^��Q�����3;OX�K�.�=04<Z��9��YM��*�N�����qƝ�Q U ˦i��d:MC����	���?.�c_�b���ɲ�:�G�SV!B�X7)M���(�Nһ-�1�Q����'�N����Iۣz��ջ��O�]`v�u��F\<G��I�������Z@A��ۆg�A+��2�0D�۞�I�4��rX�#g.M�e�� !�a�<`Q �Lq}�e�Ui�3+�l.����I���A�&HVC�6Jy��x���1�o�]��w�Xƌьh�(���#���F���k{Rt\\o �\ˢ���Wq��E�K�4M}��j�з����%�[�R�r	��ޏ�Di)tT��%q�QC�Q��u����{�_�
L5�ހ_�K��::�i���C�L31�kb��*�<�e+�b��^�Im�i��l�bCC=�&W�фR �#i��]̦2%|����4h�
�>��`*�ڦ��w�t���K<�1_��M<wœc�� ��2O>|���9v���y�ڎ���?g=�ՆFD�i>������ߒ����QRtP�ܺn����{�b�s�����I��2-%!�4W�#��vs���G��Y
;l�m�Y ���>:��\�������O�+�O:Gv��G��z��28@�����nf&TJ� ��;�����Gjf�T!��;��#��ݻu��v�id1�~�8(�&}!I'q�w���h#P��~/����	���7�h�Wy���mͶNt�c���,Ȣ��
�\���3f���2��6�-�*k���k���`�4]K���C��E�QK����=��K�	���e�w��'�Vځ������}Nc!d<�k8��v!�j��p=�O~�)u���B�?2"��H���!�!������H����y�iC�7�0��):w�0[����3�\���jW���P�%F�m?=�d�ˈ��#'e	�&�K-p�D`�0vt֪����C}>�P�zZO�8�B:V�C����Pa�X��F���#E��s��&Z��	8�.�=�m�!�m߳D���c�^�ú̟����~;u���l��V�)�7��ׇ��^Zr���-�zel´!���)�Tbζ@�պI��~å�h�F�aF��y�йG^��&��4�/D��B�}vq!���*ȊǙ���'q"!o%�Ѵ�3�k,�!!�����"��Df���}K�꒔�:~�:L�k��8`�zr'�Z�	��(����=j�R0.�&�O�iB��l>Ω��C���ds%@���b�Ev���IB�g=���>!���p�{��L�_�s8���g��u�0b4��i	C&�qM�L�ȀƳpj��T�1�LN/��hC}i���4&)9]����͹s#X>���M�'�/�D%��!�}U�s� @�����r��f�<k8z��,I�f�̃r�%���Ɖ�#�3�0��~̻}M�l;��f�ae����}�C)}��j�`����$��'D���`(: K���EI�k��{��+�fP.
�s�`�fHL�s�)������!)I9��s��Z�#x��qM�p�g<2�f���}�}���҂M�U��1G�e��DǑ:��/��t:s���cB�Ҏ�`�"���ٲ�����6��|!���ˏ�/�WF�h`"%�lf�=$b��㈧�/�F��3�%m>�9Ub�ū�
��� B��1�������ق����O�N���.r�x����xɬ�tѝ�(qUS�t�:f�Dw����%�ǄAj�yJ�ʬ��3^lcy]�S�25d�m=�.ں�ҁ3��m�8�U1�wZ��U]'�}
�����Y8oqi��iئlUc����)���2��r������ކ'	���=`*}��8cDr���5�d�`;�R���0�Nd�����_܏�r���l�����6
pB��= ȳŨ�B=��E¶���1=[��u�fT����D�2�����io�$ܩ:��c�#*P������@1x��`g�h�	F8�Or~�sp�AC����?�;�N�;�~�H��=|r]��}G�o#���g��M��Fz�N�-�V��6QK�!�85���Mɴ%�nhBC[�1 ����dt�`#��`�O��ɓ��ob�Wm�>{�pӖ�� o:��:V16���[�����ϬlX����r�g���ڜp	xx�������6GHo�;��`�ܝ�Z��$�勑�/��9��{��3!����d��PEH_a.�zzw��D �:߻OhD�����9�^G_�+N��1���F�Jƈ�-���.��VN�Cd�˳�ݼM�Z-Y����r�=�!N)��k%f�;[�PuZ��(�F89�";�@�a�459i�_���l�]�Q���:86�\~6OfkU�k���T��&l�!��Z2zt���(9�����O?��;$k��[��3+tf�i��0d���0<�}����k�J1��o����+6T��,+ս�����U�Q���&7G�fI�1 �ش+��uy��ȵ �_e�g����3RxÊ������.Ct}g,Hb��Eٜ�S�������D9!:,��?
�v(�xwF��ev�y��d.�|Aw@
�K�T�F���LO|�	n�`p?�FZ����)�M-���u�gr�M��Y$e��M�yr�w� �>tj��������������d"H�J��ks;W��c�(nvm@ـZ����w�9`���6u�F�T���9��P;�H�À��q���UǑ��qn��7���s�Q�^�(���3�c��kx_|wS��ldx������%L����Ƌ�rmn�I���rľ��L���e��"v�]$H2X�t8�%m�������k��U���~rI�T�a���M�����S�p�qT����;�M��bVUG�&k�(���WW�(YL�3��0q�ж
wܪ�>�;B�!�+�7ٌ��`�m��ay�Z�Hu>���9�%�rA`I��π�n4�]����iI�f�BՑً̓W�l�51v7�-¨�h�:3kzr�ʔ�
��*#�B^R�v�[JS\���(� nHSW��y*�b�,O�R�Ay���Ȃ�H(K����e"�_�1$2<�kPa5� O��˕��	g9Z#���tٿp�S� ��cw���G��!��V�CԤBH�{3Z��7N�O@���v�-��!�M �!D��1�[� ��)z'`^)#o��c��D�Q�����+pw������sq|5ѧ���O_�? c|��<\/ u�)�W���6iT�=%�*��6ϝGZ!��BH�E�_��NU��J
���k��]\�b}'��2��{�s.����Lo$�u��5�tN�����[Ő��T�Y.̿�_W`ꭵW�o*�ق��Jc�wp�w9яk,�۫�
+Z�.��nR�n8�����*>����%'D�*���ss�4�ҭ�{�!��x�)�R5W!^if�4��Gd�w�8q���I�n~s.DM�g���t͖�r�������~f�D��+��r���߁v�b�@�&\�y�u遏����_P/�m�諾�K����Z~�K�n�ی�l2v�pf�?z����2���ohrZ�1ff"�##����Eh������6�#C2��I��>�od���l��5ա2�-�������6<�(�RYv�$��{I�=AΖ�vE�A�$)�6���,��P��yN�S�Ku�{��I��g9-���j��D�ihW���, k���JL�x��1�$���Ru��R5ۘ��)4�]t���
/�6�,KP�'�Z%�p՚�n�d�t��Ax��Y��(���LZqq\>�_=Cb�7����)�$����p����{�Dј��xx��_Nt���zի�2xf��gfY3]ѓ��u�O�����M�V��su�`V�"��{1Y5
��c�9���UD��a����'���)7�s��!��:[�0C�/es������K���1���e7βU ��cѩΦnݔ���8�V�h��?��}�zjc$�A	(T�`��T��zB�K�=�ϓ�=��ܑ��9�P�i&GhŶIY�pd�S[b�O+����Z��p�'w�f��Y,tL��}p�H�ǥr	��;L�}������6���=Zc��NR�x���3�>D��Ze��k�牭��P��7�ާ�heX;�bJ��at�9D��`�c�X@��{�$B ��q�el��9���?k]"JX۽����G�rb�|��LՅCFf� ��0��3/��+�^��r�ԣ)�|�D:�s�v�Ge"`��� �i�g�T�����!�:~�f�q��M���Nw��8V���w���qWg����t��ܒs��+X�]��s&���<��z�ş21����t��V)�����X��$�߫�v�ʑ�d����lP:�y�0��v?0;���-o�'��2��d��� ҏ�V�[o����� ��L�/4�ɸp���CQ*�p�xh#������Vusx���R�rD��ZuI:����\h׿{�r�J�̚��/y�����D|��m����i�R(=�:RT+�KV���k�z��1���VB�(e���m4Am�%�y���X�����^�b�b�V��w���� F��#$��J�:����_C0���� i�C�Y���rm�I����`�db[Ȋb�)�ؓM|���Z������gG�U�dvʏ��}��ט��W��_1W��5�f����;8��W2ͽ�#�m���Fy�`���wB������6��O�^�� ��5k-���WK�[9�m���U^'A� /�t�I�/��R�R�j!YhQ� �W�[j�g^��U��R��!�4�'h�DnD�-�>>��ag�K��k��! 	�[���-�}	ҳ�/�c��eH��"�G:@�u���� �Ǐ��vEӛk-+�"݃�Q1�.�G�J�Z��4�Wé�Y�Y�ʮP��S����)��S�}ð��3g�y��h�R��g� NѸ�G���d��M��A�ߧ�h��ƿAu�J� ���#��9��b*a&��]{2Q-X0_U�H��f��X0��F�J����5��T�k�Q��un�}B�3?���z���G��M'�E����7zBm6K�ԧ6�B��? {f��a��s��VE�������<��8XJ���8,��Q��)��׳,0BҸ)�۴� DB��o�b4�&���9�@H��k�̥.��!L/q��H;����&(q�,m�aL��,-����]�ʦ��f��q|rX�ӎ�U�R~�`���HNZ����+M8R~�I0Nw �ȝ,�G����KP?d��RI����3����7�Ն~�v�s�W'�o��-!yf���������n�U�����$��j��4Xi
�_{�񽱫�}C��f����Q��Hۉ��S��7�:M .���[�a���ۥ8S��/��k#qp>ǭiʌiծ_/z$���ÓFE��߭�*�h�c��OB����4��*��;����P��UU,�Z����]�{���w�[�U��f�^4�T�)�xL�ڴ��Vq��=��@�r!ꆰF�m{x�*��e����#5 �TK���1^�ڸ�N�K�W�N�-�u0��K���4�돟�/T5Y4�J�ZO�Œ�e����Gl��I��kj�l)c�q���&�U�e��9Xȩ�m\<im�"K������YQ���J�U���m��U�/��J���0��3�l���w\�A���*5��}T] �`���l?>u�=8㟱��9��PՋ��`)�M�Nz��F�;�C�}-�g����,���m����(��ᶃ[ԫRt�X��'[N$l�R )zu��i�NS7U��I1
���>�)M��=�*.�#���OI,�X["�A����BX9�##�1��0��[~�t%��X�ߵ:c?e���Y��Y�.������J)8G��A�l�;�hnոr�\r�vtf�s��f��v���Q9�>T��k���(q���a�P���y|%�����9�S�	b��XI?������NI�#V�ܬA�6�@ZJN��e�9�(�jHr������R�~)g����I���cx�Z�a0����8OPEh/n��B�~��h��iSZ ��H�Oʗ�N��Ȝ��r/[u�\RMu��MW���0A6�I��=�1w}�"�",�b�BύE|p�^��I���O�B<̜I���e"=:qӁ��d��;Ē�E�$�m�̶��K��ǰ�6tx�dz��R�Q1"Ԏ��� :z�"%ʪ�A;/2�:�Q��>���3�z��n�o�1��`>�z���Tifb�$d�O�4'VMﾟ�C7f�a�wYS���H	h�"�yrr+O!z1�5+0�5[x�����>��9X�#m�;�0o�M洲vt22�I��c�D�A���)�nfg�?(�}�����P��˻Y��P�<����i����To��Dҿ~(���8����Hb��"�ڭv͠�Z��[����b���� ���?id�DzK4R��sr8��Ck��Y��Q%I�P�ezjt���d AH�o�ƞ[F��&~��PEc)8G���}g��{w"C� q��n��~�-����)�Z�A.*
�L:F�>�?�5�\mļ�u��|=�Ո�����h���E�{�*"rZ6󱐑��I�˫��޲H
�F��= � �Q?l]���d��$�B� K���SL�g��%�,�����{��3���I2������#Ka�c,��t���2�x98�	_�H�e�n�?�k5��_�8�����H�2�6�&1K֎\���G>LO�ߧ)��^��TՂ��.>�Nң�V�p�^���)y��L7')3��Jp�v� ��}��B��>_��7l��Y��EN���b�:<����wY2�&]�m4~k�Ђ)��G�� n�|�J���������o��m�Bc(~+D�<��R�z�1���Ck�c�ܕ����*I���_�U::=qd�=ˮ��Q]��{��f���r�-h�˱KքL�<E^gЇ����l��4��7�5oO.�JS�Ok	��v�L�Zd���h�h�JD�᪔v���kQVa�:eD�p�A9jld;&�Y֏���$A�H�ɖ6�߸t�{I�U�'Rzn��Ե��]��M8t�D��a��?1H�J�h�w�Z>:3jB�2&��V�Xʳ���C�O�3���N�[��Y�"r-)a�B�6?S~����α��0�aZ���3���$�9;lw41�ހ"��H"{�2^֗%Mj����Eqd��7�~�E#	���� ��:)�ޙe��лEƻW@bˌ����fh�P�����8��Q�I���]Um��Ik"K�.�6҃J����S"(j�ca9��&��+q��Io���X�=�1�}�(��s>������ :�1��k<�I��f���"� ��w�a_u���{��v�����^vnR��]r�s��{\_�AС��?�a���V�@��S�����<.�@��f�؝����:�	N;�g��/�+Y%=��6�,Q���p���d?\�<mRdr��
��2�9��9>�s��Ⱥ�耾��k���Z�_C�����#�;?V}5��3���E�����K߇����G%�W.+up�'%�z���7*��^��"�]�"�ؽ|)���`�T��̧d�9��Mc$��(k��J��>����c�u��4|�B�g2I���v�<(ٰ�2��O\��c/�8�,����4rOZ(qfY���c��5Ğz��,΂�1������`�f����U�H\$�]�_ѐ>�$���B_�~ |<��ޒ�����R�Y��Z�\�6�.�)��`������L��6���c�2���D��	f�����bLCEq˿��W�F3ӵvP:ې�
<�O���$��*K�9�{�;���aE	��>��3��؎z[3��E�4oio�����Nw6/bhV�-���"�pz��j?�;]h*��c�A�t��̵<������l�9cB��TO�Ե��¯�1����MI�۞�e��a
��������A94R��(-$��*����	�a�:
�أ��� ��/�jy�=ĵ�f*9�vpޙsR'S}6B��^Ԏw��z,�7�<U"p'�!|<c��T'<_є��@3]�#�R:v��(�B�#v����� �E��E�ex�M���-�_��~���$���`à���"���P_p�qG�r2kn�	�6^����0>�}�3�E���5q�䴋?�OX5�N��D�[y|�T8^���j�
�(��G�L"�a��^ؘG��.�H���kȠ�"�z#.w� n@>��i���L����#�?Q������H�N&*���k�����@�8g<dd��m���:�
#��!Z� ����ls�ֺQ�6Xƨ�������;�冻�g_CM�%00M����6�"�#ّy�ϟC�ѤU��򃀈v�
O�^�-�tGu�~�5J��b����1X�m)�T�Zɿ�M�;-���X��IF��\G[bnP_��I�輜���Zv���� ���B�ϖM;$�v��U�����!�7�c��PsǢK1�Mt�Wpt�}v�<��hI�i_���l�|��Gc�8��DԹ���j���v_èQ�c$h�oRMO'�~t®Ԉ�>Wgp�I��ʩ!�o՗�s؃U�\��a����2�Pz�W�#(�x�]}'���n�`���]J�(����m�>�$��ZS
2p������gm �i���$��J�p5T�=;	���Frh"��V��<�c�V9�X��ɤ��oLT�e�E��|�V��к����C���`B�q.Oo@+C����j���"zUB9��]�4�b��.B��SQ��(��=��=��C��*c����:��O|�t1���6n���V�x�{�K��E�3�vJ~(�}��N�4f�!���q�����яB=���q+�9^$������E�-�0��g�c��4Z��T/�}y�0 ��sO��_3��`@���`��,�|oV�),��0&l3�sK��̄�����<�u�c�-�(�j�H�PBI�n��̖e� A���x�n�+(��/�Nv��y�&�����<�[���v��|%��
k�7g�8em{#�И��c>mK�>�e!��x���P�%��H:b�x���j�4�3ܦ�����&�Ń�Jt�<��g�WM6��s��� �G��(�~�J�_����"n�d%�Ldϼ}R9�Y`m���`�dzyVcb�j��Ral�1�f�|L}M�c��bek a�h����lrA��`�ܠ�4�0�D��ByT�V��qI���('�P֪B��w�[�u�K_��_��@ج���q�XG���� ����E���֬�0����gAH�J��Y��<��yP1Ǩ�6Y�
L������u�&�/9���v���~��L��0$uB��H����J��r��L�8�)���f�Bu�u�:�%q���z����� �����g3���&�h��a���SH�+R�#�� ��G*rJU0t�:y�ۼY�ψ��������59�J墽&�1��H�q+���ϊ��a%]�|����E1�z*�Kko�y�~�/�* ��.���Q��9��rЖ�-y�l�fk���[��.�5�b�fj�.�D&���6Ll�C��I�oV�xiF�yy��ɣ�hQ�K4���{V��0T2���y����J�P�o�M��h�XV,R�3�g�0� �)�6�Z��9�E`�`�B�n�U8��EI���~�ҏCN�T�A�VBq�X�[� ���wz�{��>}xŮ�hf���E�ι�5t�T��n�&u.XK�*���JD��Mmo\a�D,�Z���UI�U������(M����^�(eV�� �_k���i�u[��S%)3���,O�
�w^,p��m�e���p��cZ�:iae�`|.��x̚��GY��[)T�NXE����z+��3ZшN��t+vs��e课�g��7��D\��ڮ�K��]�6�l�#��jD<&{n���G�o$}�Q0�L�}����U��7�=lJ��M�4���D�b�;�Ր]�fD��r��ý��V_Ž0 ���a�v����D�>"�Db����9F�94�:��]@ ����"��3�T �Q�!���I������j�5'���k�q.�|1���s�
k�n��ծ�C�k��}ѧ�Tlf?%�1�@I)+O�)S��PO��-Z�7c��{�-����1R�d⸹��U��J��b��)��#��gg��G��Ǽw8q-�$=>7��j�|��c]v X�&�T�ZV��~�'W�w/(������;sB�dG|�&qI?w.�H��LqX��q��P䛎2�匫=;�+��3	�.�h�S�1��q��=��^��>�;�!0j�۠�O'S��-���?�O��%�iͅ�Z��r���i�UΈS��$l*�_�k辚C�k$������|݇����73E��� �,ߵ$���k��	�ju�ŰD���Y�Q�������*ɾ�Q/�[�`��ǖy3IM,�.��aQ�x��ȊxJ�׬'{�I5��m*��Ns��1���	����t!�����I��5|I��Hڳ��lB�i
|U��㒒'\@c��)Mo��aP�˪��Ye��(�x�����v��X,���g��A�8�}��J�����F�ǄK4O�9���o}Cl��P$�s��+�vi>�������0�LHE|`�W��=0ל2�A�$�Ț�}M�F�4�o�p��Zh���B?�r�Cw�M�mo��i���J�t���oP[����y�X���0�a�Z1z�lFĪ�������æ������~��pHlX&j,�QȔݤ��"�ق�ņI��
-�A���U�ᅮ��:�=}��ܓ��G��n��v([~�їJŧ�����s����\�$l�n��ۜ�޺Qg�4���T�C��z���,��3�A@t�_�"L�&T#�
D�~(S�mD�y ٍ֟��̖x�y1���r�g�}8�MWdt�yt�=�Y�����9�e�{�5����V���|��`|>dnj�y3�W�;��uaZR�S�m��3�GD��\+�IC��j��fH��f�|G+J���A�Q��R���x?e>!�͠%}�!�R��[������j�*�I(��{r��xΜc���Fܩ~z�t�Xk��P���b��I���^r����V���!7���.�Ns�̭k�yx�0<�t��P�`Wxˮ��v��X�tF�n�g;2]Hޣ����G��`�'��~�+.����"9vo����ͯt�	��포M��=~�h�(��T�c/3E�`ʒR��D}���DnP��x�)g�� Ў�G���V�ӏ���wX���@{n�J?���!S�S98ߩUm�?�a,�#�$Ɵ�Z'��6��I�W��0�_�睔ܗ�QW'wNt0ݼ�����Ǯ�쒲9̼�m"pL%r��>	���b�E�� -�S��n�.���_ۿ��캣0G��e'���4fZ)?(�ط�������E����6Wl�Q���8A�X�H����$��)�D�6��t�?b[P���nWnٕ8�ͅP�L�����=�CMW�����1[Q0�$�bR�-�F������a��wuM�~��t1��rx#{�Dd1H�(�Y�S��9���|"���1�.=�,�
ً9��~"Ņ�no�~�m�@̋�2f�-�%d�K>��ܪ�cؑc�f�����/S��DCd%R�W��0�(���NR��{C����
��b���!T3ÂV��y��`('�L�G��e�>�ݳ��J���'�j��2�p�r_�<��S��jJR��N��Uy���ٵw=�:s�<�B(��z�i#��(��M����������O�Cd������I�څ>��`e�l=@�i2��ph�^lM����1��؏��cA���}<�O�#J'C�0p�/�X�&o;|��J?��bJ�pA�� K�Z/a�Tblɻ��f缁Tr������s����d��A<v�B��g���`è�ʨ�W�l�ʻ��h�z�Ϛ)z �B#ȍ~�Z��	6�?.���\u_�EM����ئ|^Q^��jr^��Y����ƅ�Z^ŏD;y��\����^����0���"�Sf�N՗k��L�'�׺eq(l+�fc�s��{9�G�ۑHs�����f9�������c3�6��oW�u�e�F���鰱6��o��ʑp�De2���m�E1�n/��%;o��-�_4�B�!Zr��u�
��*�#;�L����
D%W�g��znl�9�A�n�;�(��Z ���v?s�,�_?�1e=L��Hn�=Ra4����ܲɀ t��+>&�s�e�=Z�AE͈�P@2/�A�� ����_�� �b��;��w˩�7FxX�mk#�)Q�s=�g��v�	4�s�Y'z���S  �Wx^5�(b������PI��<�:�#�g�R��"z7�'�Y��g�~���s2���Zg�G��a_�b=r�]�+���SB�HUX���%��p<�X�%��Ԅ��]rQEz�j"��蓃_�>I/����<3�W�8� .�8nה��S�uW@�xR��m����6�Cj��̍���:�/�� �1n��y�9|TI�p�A����D�j{��E������.�9m�a9�{�?)�Zo��3׶YA|$�K[�l��O�RҴ"{�I��f2���d�8fs�"�wll+��؋�v?�I}-M�&9�ɨ(�㫌/����<*����� �N_��ʿ*��i��3��	UU<x�B�j�1��٤�`�O�����2�os�Ϩj�މ�~�9�!�Lڷ�5g�*��o�ٚh_��@�2�)v�g����Am=?is��� C&5(�@'G"�	��4WJo���}Vo�|[�D�<4�[�	Ob}����	&j[BEa�e�E*�<�S�'�B]哧�z���I0�v��������e�x�6�}���Wj�O�;cy��]j����v$��	j�N�~��2��$�QZX������_��1�d��2�wM�mz(��l|k(�6*���������4������AN@� ۨ�J��.*gBG���O����Z9��B�쾾�@�b�p�uc�ٵF���x����e����ć����qBC�
�V�! �T^gC��Եy��<O��{RjF������;�^ ��u���a&/��k��7�/�'P�͔An�f ��#�� �n$+��̙I��%4,}��4#9�-\Lʤ3����9v�!~����oX�q�	r��v@gN�{y��T�E�A��?������-�i�*X�ϻ[��ޖ�N���$d �6 g���N�D������A}�-N>���#�)'��=�M�4��q��m�̉�=.�~���Qlx*=#�+��,;b����"ՌFi��Gg1���Qo�<>���6�wbC���c�Hk��V�ɚi�d��5ȓ!S�F�yz[��"��͜�Mꡡ|R�3]|��QP/(nl2^<�/�cH��1#hڢX���I��:�7�� &��/� ��z	ؖGEs	������	/bʼ��3�1���#�W��:\���დY��B*"M̊���8Q���p���p�N^�0�1Å-U@k5��TZMiȌ������6�!~��Z��GQ��\�C�)�*�K�L
��
;���V�FP:�y�{WB����`��D�g�_�L����kl�
��i��H葄A�t��
,�}�R�)y�&k��GG��;1촑�hX/ɚ�<TTIX0�{�7N���UOL`����4�L%��r��{^R�^��w��o�K��6{in�Ј�%�Y��5�V�ӕK;G�0P��ar�]�}۷�E|�
���~03����-���/�4����k+�@ {x�3��f���1���Q�K�/��o�6jX�s�N��KJ�#~S�� � /��O������6�Nn���Kg�R Ɗ�`uey���%V���8��ӟ��A#�j�,���z&�#J��ր�� �*����߈w����e:O s-͖��kC*xXq���4�0_h��r͜����HzQ���v���޻�; �5Y��u�9S5��QD�PSj���'r*���2}w�M�$a�^���{z1Mz`p���1}]�.}6�Cs�p����X�b�a eX��,i��kG�˭��<N>��_�h�k|�LՆc��}U�k�Op�DG������#jީ���9ŪY*��`z�vD����a�1�!�yRc���S�.18,���#� �F&�k�+y�cI=V�O�ν]��S+<IT�8�}F�����u����:w���|��P��ګ
,򟠐��n�	�8>IC�jr �����2t;��_���� �� �������>�Υ��;��%�{m"7��m�;:D"[���<�Dk����{=��b
�Ja�T���~�.��H�;o�����SȚ=,������`|�GO��(�
d���n�\����!7�ŉ�� �����x�22�+��|5��y� v�]�!J����۲"�v�ؾ���K�կ��hB��^�����;NUN\ ��VׯW���
e���F���
�>p��O�������!\�D85lq�9���}\���b������k�A�js<_B���r��#�1���y$�����~7����ʵ@�Od?rwZ�M���P���m�Q�s���'����Y�^y��7( S=����k!�b����r�#�4��2��bpC��R+���I��F�x̿2y�:3n\%���J���疻Y7V��g�$ޑ��u
���ZU����sh�=g��ەy,�I^-�=������}�����Ic�ϛC��'�v���i!6o��}x�U_�������ҟ4�-Vt~3��D��YjUx�f�
�馐��P.�!ĝ�����C�'Vl�p\����Du�� f3`���o^8�l/	���*�~3R"I`~��9S�fJ8dP����nK�|ls��t��*��g���7Z~d���)}2�پU�Ⱦ>�u�R����CG�lі��fR<n xA�����Ŏ �<��ʆ\U:�4B(���Y-�`Ld�)M.�)��}&2��s�$a	�%zÆ��7�&�>�u�t�݊;1�mVކ��M(�ŵ���PYmШ!�y�}ἥh�N϶������g�'�~���/�.o.�O��' �@���B[%^�-��A���;T�i��I�p�[_΋I�M�Z�1P=����0�+c
��7�O�J��^�6)�sB/�Rв�cu�o�]"�WG�js���i�v��������r�\�A�oЉ#��8�/�ErO��<�o}�(���v�k�E�\����ġ�I��x@�%P/*� ��y� 9gk�K�q�g�c��o|N����ȳ*�L�H�b�=E@SFtot6���+����.�#4�5�x9�m�$^[0�:�:N6��Ok��2Rڼk���I���b�Ww�g�@���1s
�ZZ�J2S:�1̝(|.���")|��Q6��#!���|���Ɏx������7�]��^c����I.�U�J�cT�i�hz[�$�C���`R���+�r��W���m��d7�K"��c�4�#o���ۛ�L�Ae>U�l	s��5�E���/� J���U����=�Xh.� �z��+�B��f��8m#��Ufp'yp0�8P���_��XM<�l� �>��ax��}���������L���6���rfD�C�Gw��9�U���w�;'xg*�=��t{zJ[y���m�`�I+P?m�]^����=�^�C��P8 ��b\����D��k+�꫞�I�ڹ-�*��V6�7����U*�OF�a�ݏfM���/GV ,��EX
C��"���oV`|o���ɗ�ORG'r�5ڰ|�d�i�]�:���fH%_��g�#~��A7���׈`U���y����&�7�F;�|�
�s�=�+c7��Uu�Jt�1�W6E�	�6r�h\�4�@=��� Ú?���oOݱ���c�����<8�mweI��Y��O<���ïဝ選W���&#[��!��6�ҏ����U9l���{��v�B�Os�)���}1mM=(VbU1��'*����f1m7�t��[Z��z�_ε��JĽ�JL��f���Y�f57��4�ey�F�C��к�^���_��l3��yf�\��s�܂>����Ꮖ��K��^C�����b���Q�@�a�G��;sO_����-�Ra��!����D���ۙ״�����v�CA��1Ӟjd�+�o�N��'���:�
�O�mϸ����R�q��!�#2�z��D�Xd�hLA�I*����6�;�%[��Eԡ����x�S����*|��Wԇ��<K�!���s_���nPl4z�?�g'i�����A����ӵ���QC5y�ѻ\���G�wk��;���� џg�`��/v$*��!�ή!ш/��Y�e�6&[�Ip^jA��=s�!�91�Ub��/���~�/�::��fsX/�	dG�뻖=^���X}h�8|Bmns�v@ʵq��AE���ۿ2�Je)����cQH}+&����ݶ�d��V Yk�VIA4⾊��K}�����W��<���n�c��2I�ha@x$i�
�1�$S�`����l��g`�2�$9M���hX�I��}�n4s�v���.�qk��g*[�#���?����!���������Sr�E���B�~�#Xv$��ėԾZq{,4��T ��>]��FP���}t�#x���o��Y#��5P���p�!�[25����K�hjL��~v!���_ZR�a�k�������ar�>�B�MwȬ}�� =MP&0��Zc�[�[�������J��k
@�~ל?.�g���� ���X���n܈�	��}�я������0�Jf��$��Ş��"��{5�b������+��2�!c4�D_Zk(K��wCE>�����~h=�����_��^8>!v�`5����ƹZ[~�v0mk<[��Ԟ�Ħ�Ӗ^�aKs��f��5�>e���2�K�R$�ё)��Ld�dp����nxծ�Wg��=�\����N�n�X��'��X�<��(²�<������ʁU����[��;|/3���lA(`�;m������c"��J��6d����_�� 'y"S���sx��&^� -m0��!��˭���\��M������;�{8�#�G�"�:}��x��4���Y{�Ϯ��?������W�m�JR8��P~I�ykL�G��������ni�4�.6�gI��E"W���U�b��C��zXٸ'��\��H��#�����|��X���bu��8ha��=�!���E�|6�}?o@;�pS�CB���U�R3-�Y�L���� �P�͵�J.��&4q������2���+�_v�8�؈�� ��� "w�0%TŤ��<s����\-�%p{p|��w��ƅXd�O2��Cᒼz,d�ۜ�ᦣ����(��N���Њ���S�63DK��j����.6^!fT��M+���x}O4倶�X������E�j��@�F�<��《Q��㬘�����=�_��(�m��7�A�`P��O�F��Q����������F3��rf\v��c#���U@OT��FUa��ko�D�;6ȔyW�}��/��ʜ!��l��^���;
u���p��2ʰ���~����2����DuF!.��M��態��q��'+�l�@�
A�F:k�}`���|����؅�4�1(��J��D�� *�D֛�d6�/ح��8*�1e���D��s�k�т㭣b�5�?:��]�����<�,nr����X?k�ݵ����a��RT��A{����/)�3�Ĭ[��yA�z`�IQ7ܕ6���%o.��������m^c���4��xE(�F~a��t���.v��u�;����B��Y��Id&mPV����I�$ѹ�f�`Ov�@E�:��h���nz�!�&�����q�*�����w^��������q'T�.�����z��dMjk��	kv
m�"f���Ea�Tl�L� ��Ncs�	F+�uL�ّ�+���������`ri2g�n����G���}�e����`Y��·�rʼ�f�>��M�AW�+�����rZ  �.^�٠���:z_��Ήj���*i������"��j03;�"/"� ��S���!���W�!�Ѵ�zJΙ��1��@b|�c�R�<Z��=�>��KX�	0�I�nD�:�e~D��ʺ�H�����G�T߭_u�v��24��Eo��s ��(,Fjj��"A	m
�þ�r9����R���W�Zy��&��� �PM����|wpf����6���7�uJT߫�Ad��C�#V
��E �!�`�S�b(�ák����fP}��ڔ+Z6��a�ءV|a�C�!�º��B�o���������y͙س����GЊu+��pi�n+3�:�l"�ϗ}��U�q������Su�x�"a8�ν w�[4�%��-RUL7ۯyށǁ a����I�P�W������D�����{�?y�8��,����YL �B�G��AS�(=�)�+Ag��`�M5 ��4'[���J��䓆#�FDa�@��ה��5p���9&�mOʮ;��Fr�l! �^�:�
�iF@�T8�,�F�e����_��n���o_�.<�	�.��tk��̽���{�Z0��îG���|9x������gFJ�56�&'�ߝ�vL��-�18�S���͏H���]��٩v��D?�Pp���P��Yδ</��Nꑾ^A�):7fJ�;5�+jF	��͵��Ձ�}*�#V�����H�U�Y���D]�X� W��	*px�s��bJ�s���0���^P�1;��2��������k���~���IԤ_)��O��cX�nD^�5BKt����h2A�3?�{(k�ϙcԙ_2��!���!n�+=��]���Z�_�12����a^ �͜s������I����*�K���s�� #X�B��SM=�	��(o�i�(9F;5��( 1�#�Z�����L��7L��͇�6hG��:o��{�Fc;rN�g]��ƞB�V���Ͼgv�Ȁg򚋹P'H��!��s�Í���l��4>I×wt�v��aչ�T'$��zB'Ja7;�n���/���w? �Z'%t1B�F��cF}����VG����Tu 狱��5Axa��Y/��4�?;�&�:�_��3��\bHuZ�U�Hفr��f?��KA~�m��Jߥ�q*���G@�c���8n��X�_�ҡ"�#$��ܿ�<a̋��3UBxʴd6+���}:�\^)���/
z�:#��;��J�����!��6A+i�Ij`]��b�eT�(����3��ӷ܁/�f�dx�S� �g<�:���N���9[G�C�_8���<�����g\ᢚG�Y>fHa竮�VG��7Q&N{��O5���[�ĚS������������3˽�BW�WK��j�/����\�r�C��N���3;{M	�i=��o17�{�/��-�qX��M@�r+������VRs6J:��/1��&+�����g�a���|]�Uxq�l��} ���rA��������*���aWh�<��_�:��E��rNl���ph���~n�z����0��O�^};}�#��H��衧�ѵt�Ծ�X��&�??�Y@�����̬ka�{χ�qQQ�/b����j4��8*�;@�CQ?i�Um�و��9�誛��ª�<4a8/XA���ap�rNo	�n�3��ik�j0+F���̮[<����DȻ�&��㑘ϥ������rp��'���9hB����k+Z�>��H�c�����2g�q��)�u���U@s�)��K�^�"�ο��D�zs+0��>�1<`�K'���!��%<�f9sV�[��Z�J鍸g�A�ǰ��Qﾹ��)����y��%�s�s%#��� gͅ�M��q�6_	��d����f�t?��������P(ܐ��x�!.P�_ˆ���P�p�C�\D��H�Ex:n�@��\|Cr�g����!{� ��.�m���>�x�7�,I\4��x��Tn1YNP8���f���%�����UÝlŎXf6�>mb��@S�QN���w�շ���b�з���vP܂�/�cq�<n�qhEAG1�!J��ѦH<����!��,�5��������v�e70n��L?N����@v�!����
���橈%�?������]�:mz��5���n�\���1��
�n7b���A��u�a_��G�L<�j} �,!>�t���,�P����7�����:�D72�8=9��-����,m��axR0���p����x���n�&9��	\F	5��t���R���f��}8��9��j��(��(�/����k��ɓ��D���Z0���n��/}�쪶1�����������Kڲ>W:�W��.9�!Yd;菉:�U5F�&�G� ֒&�Җ�VۀP�N/�-*�9��ґ��k*Sc��v"l3Bˁ�p'����_��梦0d+��� z����<��R�~+���07<�1�6�V��i.o;�L�q�nI>�]N�]�`��/�u*�E��ݿ����w�?�M�%��9L;�\�U��"�.�u98>%���CB�)<	�\R8X|�Et�(��L���aY끺��vt�&t�S;�������I�ڽʐ�b��o���6gXyȭN���������g��:�B�� �&鹣N+.�|�DRx
_��&e��a��⭭$>����~��֪eJ��o�<b�ƛ^�A/�XT+V7d�;����-�A��Gf�u�C�a��_	�s��Zx�ZL�I�g�����U9�jŘ�f���V�!���� ce����k,�Rw�M�,����*�%;p�����F�:8�{����@ۥ�������.���jS�d�"ֳ�)ة*�����l�V.�I)}�#���+@��A��>��:Vv�,3���-���-���>l�9��3��'��>x�(A�g����H��~�Kq����sO���<XKO�F�JӠ�8��6�P3|��X�@�TZr�˫��y֡��TIc%ς#}������1�"����|C'6���9XƈAn���/b�}?��h;�ȧ����窚�-m
�U�vN'����͢7��Z��t"f`���>;�̆怦���k��A<��A��	�t�$��g]Y�8������f����nj�$�-�"��ײ�-�A����0�g��{0B�d����]Fd�{2��f��پ���޲h����pI���@�G �ME#�e8�y�����\\m6i^��G'�9�s ��1�C^��/�H��/�Yӹ�:��CzSe$��2Q�R��UD����q����~C��g\��=x)�	��(C�� ��O����d���e6��jSi�oY֒�j�FZ�B��5��_m�������LŵP�	^�t�߷Ԡ���q*��k�4�)� 8�r��:=��I5dT����.��Y��t`<��s^�e	�*˧&F�|z$pT���2oL"+:�[�t�jل/y\ YS�Bf����.�F^;��e����m�tW��G�$��`�L;�3{I���1L)ю��>`�-Z��3�O���Ѣ�~69��٠�3��m���:�&��~����㡕�RB)��L��0(���w�y*������GX~��l*k��
-?!����������"X�6f�6c���\Φyg�LOF'��O��_ӛ^�p����:R�rbB������XE�
>�,�ԉ1�PV�By�i� S�J�� ˁ��	/�\tP�(a&�?��/�oA΃��T�+����)�Թ�4,ъz�*��������.j���*�雕��D*DI�+����
�&�F%-\���&�_5F��+�^�zo�ݐ̼<D
��,=�j/S+!Q4�J�$}��T
���՗�M�M�l�u�`����m�e��,�^��Vd1.p�ⵟ9�#
B��b&j�Z��$���u��4�@Uv͝�S<���`�i=�
�Qx+ů�6��P�Z�P|��u+.1*LZ5H��)�R*z�� �qyf	s�E
������δ�S��@&��x�D`4�����V~(D�Sx���I7�gl�}�g�FT��>��p=�Lը��(e9��W�ǜKJ��Fp�Ѱ*��KK��n���d�!~^>�V"w
�?
��UI�`�Ż�N��Є�pg�YGCϯY�s)I�.��?�!`&sG�:>.����Ө���HU��Wڲ��@8�,�+�Uq-���P��۫�G�/fR����vFXƘ���-J����� 1���a9�,ٯ*߇?͕�ɋ|���45��9�/#D������@��3�Mhͩ��jW�m�����̮��>P�,�A���˕㝅��}�4���1���h�+��K�[G(�LNo����A�N[����Wi�Q�ST�}��)��_�"˝����jĆ���{^�ύ��[�S�P+��C��-�^��R�>L���o(����;����vG��N��t49S��<�U�j����T�ndB�8�.UsJ��	���Y��|Ŵ�UB��ޘZ^V�J�jOi�v60��jB�-e���	g���H	�o"��������,����><d�v��_��s��c��ib��G2�	�z��z�+[//Lݔ��&������#w�l$`�W�����ڷ���g�Ք�9���0��}-#O�Ri�[�>t�y*x°�nΛ�c�E��gC���.>�'��n�xɻ��b�-�n��Z�ӽ�J�oNH���Y������\>)�_+]c謇�&k"�}R���&S�~��/����t���<����k�Z.F�}g�%�,�l>"z��5b���Ʒ*!hD,�P��%.���сE�19¬�������)�o���ǁ��������F�Z�
��)�}R���p�	�&L>]ۤJ<�:���U�Y�>��S����@���_�t+�p�ʯ�v��O��7^���'��5=�K \�ŕ(����}�z�D@�'9/��J��9 q>��??8xR�H���<���MCۃ� ^4B0���0GX@?��.;wV�|c�h�����R�~t1\��݇�7�g{��6�M�u�!�:�Chf_��2d]o���yO�e���F0"�JA�KsӇU���ɑoSW������3DC��&����`7_C��R���(��d�[�\j�T��q%��U��ĎO�}���*/� e��w����������2g9 ����I.���]���/�� 0ܰ��'h7����A7��u����Q���>��Ό�$��-�%�	l?]��^u1�ˀ:Gg��>(cT���W�[�!Գy���ꪇ�����v�)��&�U?r�D�l0�E`~�H�a[Z�xf�q���l�@ܞ���'���;$�Ǟd�֝���f�b)BY}�]�CQ�� C�g���E{���:t)&��n|�
��Z(���t�cY�w?H���,�]���=�vcg�����;�1~�=Qθز��"�Δ��5�פ$��]\'�QkG.���)�T/�G`;����S�rĊ��`p�#����#ˏ��*j�$_���+	����%y�8�"���0�89">g��fO8>嚫\�	c�P��(}E�踩��V)E�fF䗥XvV��M��VsN�P:$'�aT�S$���x3z���
kE!��C�i����ܤz�pȶ3D�=�-ß����JT�1AuN�o�`vf��i=�Rt,I��4��'厭gE��'�nK������&�R�|d�Ob���S�]\e]o�#�(t�a��`�]�V^����I�x�S�*_�k��	�Z�[_�pwd��^����:�����x��Z�gזa�gZ\�f9�@��d��xC������Mz���=�$`2�D��#.R�䏕k~#M����֍���%��W����K���zV�`8��p�]�4��Up�3-y�F�~�nҮ��~^�`Iތ=�C|)w��.2�\U1���{`I��i� �E|ZPx��0&����ᘊm�8��Q�X��s*����3� �V
l���e����>[�g��2�aih�ױ`yeG������P�4k�@�urr$�H9��������o��K�Җ>O���j?��M��{U��m�[� l�7����+X���Y�&��n�fD��V�į�Kш7�p��Ɓ�����2u�����d��s<��Qd-����v=����.P���G�γ�E���"ҧ�V�[f��t����Q����w#�~LɥE�r	�C��S���)��G��$}��:�[>��T�Ŕ#e��_x# �;KC�M�d�u���(eod�b�0q��ƍ�
��;N}G,�N�����	]�(�Ќl�Z1��{�O�߈�Z���N��DX��d<�\R]�K�sP��C�1��`���	x�ڎC������⬕��dU�ޢ�]L���|�o�ly�wXëG`Dd.ø�c��غ�9��(��(�}�$`�*o��Y��]6(����ɗ�X��BgO��vX�<ߌ.a_]���[dg"����6}�u����;k;�K���b�6~����ͬ}�	�l���(p���Z�.���Q�e؄z���N�gt�'H�"��e{��Kd�|��.���ҩs!^��i%�6���:�`�+�P{s��ܧ����ͨL"�[Lp�FP��P#�E��R$�}��^����^����3'~s=��8�I\�q֨��L��}���
��+�k19F�YS;?���C3d����<�c�B%W4�����
�/� 'Rs��۩D+Ԝ��=�>�Үw�9�.�V2���g�<UK[d�xh�Y1r뾁Kɔe�"�����d}R[%�)*m���|%Q��\˯ݍ%�`���d�	�`!
0�h&d��(3��Ru��%�؜��pHs �p� �f���n��N�y�]���@ZL���MC���"&s>��<�q��vu�(�0���I���|T�����&m��[8�c�U�Lt�EvHj+��e+���.R2S�5�[�l���+���e�}�g��4)g�f�@A��Z�����:�7��&���h�ٙi��Sг�<RRt%�z c��!���W5��l<Ƀ�2�)=��i@��³x��&�*�ܨ���y�_�;A9�%�M��� ��j�!��E����a�T�xR�����R
SU�C�>$�P_�B ����@�ջ�I�7�X	D�"?ӣ.u��Do\����]��Vܴ
d�vO�C~�w�g?ן�r��&n�K�Ip�����wI���o(��?|� 3���c_����+խ�jG���/g٫����H?(�p�d�
�����%&��(�=����~ת�}��8@a�b G�:d�s���WI�@�h��0h�Iu���\���`Pۦ��	JJ��J�D��������n-L�K)O0�m��HtUN3�����GU�������x쒊�;^2���9�s:-�+82mYj#':���jxeIB�Dصws�0���Gm�P� f�<�g'��hDH~���00��+�5�'����8VW�y�^?�G�Z����A��T�8	4�"������w���T�Su����
�%����B���喙�n��W>��3kBQ�IsY�[��>,��̱-סe�c=�2��֠�+`����m%T�Iz�^Z�L�VxW"�5�g��a��Y��#��5
F6�$�7�Q�����iMF��{�� K�����q�.���ّ���V�/�����v"|݌V��N�%.��u�`?�*+�~n�\�Icg����립>�r�4�n� Glk�H	����z��k�$V�i�K�G��s׭ �� r��}��~�*�v�E$q���^� M�(�s�m�zD4��#�9�>�>cR�t�}<�����it��:��E{�dOy����D�dɼ�G�B���:�����P�U��# ���W�/Q�f���(�Z�uT��OI�q�b[�L�F2������f��ՋK�@}��,�b���M�3��ƭQ��p����A�<d.,�Z�pV��ֹ�!��1��^��{U�7�f�컽5�G��^�G�>����$Q3����s)&t��ƺV�8\���?��?�@Q��)4��v*��S��k��C�ɡ��q)��g�h	J:}�nn	���Y؂�G���.���Ŧ_b�W�2>��\�!}�9KQ�N>�Y�4�/)L|筼������V"����਍�\pɇ I����OC�V�L�������@�4���@r�] �as��ha�)�WkΎc�w�M˨��ͭ�a�]X8�����"���(B�C�@,�"�'�G/J�է���i{mM�5a%G�%�fV~,7�-��,/���4�#X1�o|���f��<��T��!�M�u �e�a3���<�����f�[��u9��SZ��#�(�~/�Qw���M����M�Қ�����t����q'��AN|��gXcb䕞2l~y(�afEſ7�{�.y[it���Ń����,��s��l�]���ٻ��I`�Gt������"`2�B�Ɛߔ��.��yBI܁��3��c���b�I���Iؽ��,I�.�.�tY��	���ѷl��ˉ�(����ٮ��f�>�"�B���T�x�al�F�?�J���?�q)�Q�)}�y�+�C�ޑ��<y:*�?���q��ag����(��b�� sb���h�X�I��K��Z�}^/�nD�l��an�n)��o���>�	ч[�6A߆���y��T�ks���\S|��J����Ŧ��M^ٯ<�OC���;�q�?�B���)]A�a�]���ZQ����s���Щ�U�������3�е ��n��Z`��$�I��7HJs���E������T[6��{���s�I+�3V��6��-�܅�JM�u<2=1���:O��{K�-��n0V��g!������\�^̕G���z�&��/w��:T��4o�S5��V���	|��k��Ɂ�1�L�����4n��W#w����81���g�5�$v�k�2�4�5i�O��:�̌o��h��`���"�C3�tέ �_\��vi�~���]�4er4��b�AP��'�Y�YC�L���<�)�v�x v?�_���6ȍ�5�IĲ��g���l��7'|����نT`�L�&��b��=��~I$,������y7�_�0!�-f������h)�-��v�w��8]��8d�j͵�Tt!鎓��a���iW�����D�t	�-6u���ر��O}������3B� 5Ø�ń��=ڗ8'�
��X��(�<��9�_c��Z�7/�zMI_���_�������8o
p{��'@A�����B���3{�>�L��S��-@��1yT�ZT�7٫���*C����@��G��Ĭ1#Uz9��ϥׁ�]k�w��KU�4$��  �����{ӘU�	Z��$�T��"U�R�l��A�>�D��Y�9vj!%l)�&�M�X��E���W<=��y�y6�lH$��årz�o_�4��$��h�]��uyF�<��]lb��@J��������&.Ľb/�J�BC�����/�R��Z�C�=P;���{c�D� �9��<���i_�wۋH��\����I�a���Fkn�h��Q&zf�9�T�����$"W!��~I�G��EX�YH��0����>eހ_�#��Q6��a�\�	h�du�n��0s�(
殏/q%io��i��Zl}s�����C���^G*�����6I��H�Ws�)�Q�.�WwK��Ƃt��.�֗�e��"��TןE��t�h����be�n9V���J�.��٬�0v�^��]kSv�5�j�ߍ��<��\�<�^W��7��&O	՚�%舂�t)3�N�ۃe��Z�;�F�!���c����p�x	Jv�ÌcLo�f�~����M)*^��L<;����X�$$��9���tTt�e}�j�J��ww�X�����-�i����,	N�wh,^Z��QSnYX�d���F����vw�x�,&��Z�����<��вaۘ�ˉ"�3sSym��m 3&���l�#�rUf������U8"�V�7��QM��n�fJ��Ov� Nۣ7��(#�EJ~��v�/%�D~��Kۅ�|����q�M�Ă���4W�3����}�����Xl�9c�g�j��H��-m��B��ӏϕ�Gmˍ�I�+�k��a���i�ag�ߠEG��,rs0P���ܤ�n/�m�����1n�G�}�����z~MlW�Q6�^vZH�Y.�p�8Ύ��<E�z����(��׾Mk� �MN.�ӧ���N@�#�Bt8㐐+"wqC����3|��]С�I����ALT���څ^c���=�6@i���BRՈ�M�.O��K�޶�n{� ��ٱ�GS��'�v��4��K������T4�����K��z�UI���V�*[eS����DW�\z�g�iL�Bq��y�Ӥ�D��6!%��a\�^?~m(�H3��A�!�_䵖B1�l둦�_��]׷�$�����W�q�p6'c� ���y1 b���y]��xQܠ������r�Nk���%{��_���;�Ǫ>�N����S�K3yoP�Ȫ��T.�aܖ���#8��%{�{�5.�C�O:������R/u����%\��%�=9�e��-��\S�\Q{y��gW��>���ׇ��N������J@H˴�6�=���'��K�6`��I�3/��>�d�DD��)K~/u$!��SXR�So�}����c��i����ݷӥ���s"rNs	���47�	9E���J�qvN`�(W�f�(��4IT��w��}���K�c�Z�l�:tl/�ڹý���TR'�W�����lg6�C�c喾���7��R���Q}�����m'�7�F���K�c����S�X|��gTЄ��o�$r0��\^7��K�i�O���72� ��>�-�c�7���wW��滅��~̶��H��i����>�Y_�rc�q/��?^�7�/��?7��DCxF+�!��;�h'潻��G�1�k(4h_��&�f���_�^�|��Y��j�n���?��
&��vrnʧH���2�sI�{撒�FJ����E}��}���9p�?�b�,hM�,�|bm[q=ޓ�Xb��B��Ru>1�j��<�\KqR���8�G}�Y7f1�a L�_?����b���D�!�Þk���f"P�Y �%��������
�Y���@͘���̊"�Xd�	��b�@'�vK�[e�5��ڐNS_�b��e����jN���/�e@�2ܒv�h��=���M�R;�;1�^6G+��_ >Ck_� B�؞�\ {{L�C���V�
�Du�Zq��Dɿs�ᴆM���K$X88�c���>:f��f����K���|I�p�A5<ǜ���>�$���ت פ�^0��5� GJ���l��k����'�A���|:k7�~�����9��S�d�';�L���c�1������n�Zl)�<֝I8�U���-��L�@Bo�v/�(�B?��huׄ��[��(���=��GC�b}�������m%'b��R��D�4%���//�����⃐Ar̷o㯃��ۦ��,�	BJ������qA5��1Q����L��LC���Qh4\2���z�;V��;q�	«����5dڰ�`B��&�2~ƴ�Փ
��d�6��f�QZ�~�4;���v12����<(5�;G�<�-���D�'MT֪`)�F�sld�.9��s}+��R�@�'oEV��o�c�ӝ�x̒+Ј��ԁ�!�y��62#�˾�~�O���T���C.iظ�!�=�f�ޡw^�i⁗��$�<��I�ű��<<�x�����|1���\����������(�l�G�s)�,�dD�9��2���y �πq� df�U�!^E����6ӭ�)�����[���t��ʝ��Hhe���v�%z�#q��O�����	on�s��k���d=��v��V�Cb�C���GX���Y����X+:�F���0h�tM��oC�6���`�Q������;��;��)#��ㄼh�2���'�%g��js�}��PM��	b�`��P9�p�r����tM�J��|E�TȞ*@`M��D�N�<������f@�a�7ߠ���~ל�]0l�PU9_CC������ .�����.+�4�������2�.�gn�i)��/P��d����؇�\I��2KΏ����e],�E���;���+ܛNA���-�ʯ&�B#�r8�T����>͒M�I�������ǲ ��#�����o|\�Y���O��&o��� ��nI)��AG�KdA|�?ǡŤu̔~�N��%��|sǛN ށ�&a��ܣv�5܎RL�Y���G�od����I(�PI�S��ѵ�B�u&�h?�$��{~!K�*�Y#K�%%�_[�=�-hi�I����"ЮAî� R�\���w����T��
6������@"�k�4>3��逵,Q�����!�����"B���ח�N& t�oz<�l���I�,$�	8!Wk��rW��0���>�g�(����0E�:*R�굯>�͘�/«�T\��ۡ�aŅ�c���^��(Y�v���:��-�sJo?%.>r}e�� �*CxB_T�����|�c�Ub}�O���ɺ��w���@eS)�*w�..�_������!۲�U��n�텎,Oz��/6!�˄zRtŻC�M��ni�]oK�y%(^�X�`i��B^���b���E�f���y�F�0�_U ��je�� ��fUv,��O��mэ�����F��!=�6��$��9�EZ���ێXmhB�F!�̒^���sd��[�=ICE�kw��f�N�3���T-9硍+�<��]Y�v�����YFd�}��&`�f�օ9T���j7�kX��9ء���Х�*l�ys
!�ǵ���L��bL�î��@e�<�б>�L��10a���C��3�M����g&G$�3��`/���&*i� �����rP���	O�h���I(#���� �Z'�o��	��($B���D��V���h63�&����WӘ@��rI��sg�*R�%C�W-[��m�>1��Nw�񑕗���QnB�qC����b��^Z�X�ִ����vĊfy�(�~Dz�(�c��u2n_]l�J�9����)�����X8=|�I�Ҋ��8c�4�:��\�uXZܔ�������D�^�0ua���0�Gr�v7�Y!�Ke�d���A�홷әºaM�:��)jȍNȫL{'R�
��A�F+�i�N�eӭ���wa�T�n����K����MZ�H���b���䬋L���n²��E��n0+ �m2�ھ��Dmfx7åУҭ�9;}t=����V���S�]��@���R�_���zBw��
��5���I�D������Ĵ ֋,��%`�� <��+(Ό��#	��E*�2��@�"64�Fq��XwVzB�X��lР�N��]����`��i��;�����SP����|z�`V�A�t����^�	�3���d�P�f�@{ʝ����;�: {kF^��T9��8&�IH�:�D���
	M1�����-P10&<D�~���3N)�������弻�6t���1W�ZDz�]�0��ͦ�y.���RU�K��1Ww-���Iwg.G�Ͻ׶��j���Λ0H����Hc��k���a.��S>�#�%��/�K��Bp�&~~��RQ�1N"O,��UoL>����ra:�i��z�;p�Q"!�{:��.�}�B.�c��>�F�?�����B�`XkvKڄ�KbU	�F��Ks} �;��I��.�c�m~��%-?��f��Ğd-�m�P�O��BY{%���q;�В|��K�Dj	�MR��Z6V�O/e�*�#o
n¤���ҵ�"��q��x���� �
'���JL�b�2DB(�L���l���~0�F�S��|�S(�?�*���*�L�S��Ð���횑/g�/}7K�;ݫ�͈Bm��5�3�Aϯ__�N���i�o��z(��Iv,�دu�I������N�U��U���u�3�qz��8�k�@�+�4���Pa���E9,;;��P�L@YQB��{}nH�*T���}��}!n?@�ˢ!l�E|�%�)�H�ջ�%��G�����c��j��.?
�mu�,p�n#��eW;Z!���M\�*#лU�]���3�3酭x�b��e?da��|��9foǋ�����UC_x��I����ڱ2A�С�s@� ��5��5���l>7�/:�be_҆+X���e�E�w��đ��Ei�0�:�lSۅ�L��He�ݫꁼ�f��f�������ssB=�L֡u�e<�s-� ~g��؈5 D(��o��#���[Ӓ�9��a�lk4�p��y�XRv�E�OD�j,�G�xݏ�ܛ�r�ڙtG��]��G�����o�GK��m/}���d������ b�7Þ�yC���f@ľmlūݣH��v��E�R3�K�S��=B2˰�'8dPS�tU�i�'�$E��@���ʧQO	t�3�P!���)i�IXc*��	�g,]f�]�\L�g�2*���|z0|e��ja�D�$�:2m��_��n6#�GS���R.��ƴ�?m���y`���8���y���[��?-�\���6��L"p sґ��-d��`���rT�#܍�ۢv#�Br�($�Z琀~� �ަ.���u2$_rϋ����Un�	�Ns-��WL�3{h�o���"��9���j�h����Zy�ԏ��s�9�Z�I�	�a�։r��8�d��W�bB��x�y�<��U�>����F��\@5Y��o��yg{��y{�EF&��,�&�� 1$O�,N� h��,����i����6�ׄ��B�71�5���/�@�I%2�,d��C��Y������y�*��L#_i� �������e=%F�ʝ�KdZ����]?������.1�x�La���!����4�!�i�	�6C������s���ѹ^�8ȡ�[�d~7�]�E�c�d�j^o��蝘�ɃLM9s�I�7 �(�I���m[8>h�%y�5�|�i�_{��6v�@����#�Ě8���[�[��gh�vՔ&�iL�bkh�b��r��q��dx�h��$6�_�X����aoE����)q`�ED�~�$V��a�sR�b��_Y��d:-�6M��ˡ�i6#�A7��@���"RJu8\���-7<m[� b<�`am���D� 1T:�j,zn�h%����@&�{·d�ŜN������Į+3QNX���3��:���n���/T�)0�Q�2���^S��`�p�]���~�2���̓I���Uo(RJ�&$����*�ţֲ��)萁Jx��P������;r��M� n�L�6p��K�x�6�>��#��gH�.�)�E��w���0�u�O�o�cW퓒:�2ީ�L Od�q�n,��_pR���*Z������l�fC;������PجY���Yܠ�����q@6����$uS�m0ý��F*���O4&��2)��d'��Q�m���Uڝᳰ�|@u��� ��G��������<�� 8��Zj�[�����(Uϒ�b�Fw�o��#��E�S*K�+�9�%^���i�S_Y�i��F����}ɽT����)�lB<�V��p��o_f��l��w�	��NH��qJj�D��ۭ$������Gۼ�����:���Q=�������#H}�>j�'<FI�Q�e%ʏiE�v��^R���EQ��� �+;�_*1�g'���d]O��߆�v�=�Z@l�'ҞU���u�v�	#��P�*Z�0A�R�X�3�pћ�-;Kzf������_`;G�VQ�}F���T뺺>V�ϒ���nP��2����޿.L͑J�7��~���L�$���MPVB}8�{�L�JΆpVR7Ч�X(��45�����0�8 ����f�`��W\��j}��#z�wC��!!l#�f�vM��ߎ�B�u:m����c7 ����֏A?`�Ô�cB��t�1��C��М*��� ���YD�HN�@�3+�B�%ib���O8ax �o_��y
��.��4]"�ʠ[1I w���v�gBj;��q8��WR��HԊ��Kz��ɢ4��j-�A� �L�1pfeC�r�H'��08�܄,�|�r9�Z�>"ޝM��ѝ�t�,�&��e��J.�Y�]�	�rз��F2���_ꬃ6����C�(�­
C��H�����w�v��a�QU��UA���8�>A/9�G0�`�8:�ۜE3׸#�6���MH�߇_qH�v�v`ء^��-(���@�/ 덐�;6-Nb�ı�
|�t$�1��C�i"cS�J
ðLN�},mw�L�Яu��!�����Q	�l�g*�'� $C���y)��B\��P�s�q)����%�&o���R ��؉�G�G3�JUZ�+�ZO���s#Sw� ��3*it{�6|�3?<c �Es�5�<c���	��z���m���e��@�[����pٛ���~%}(z�1��5��pR'#�KK@�O�
������C�Y4�Ft����^�\?ӧ�-��j��ᕝ��}��u���[MA����*�J��#�_,-)�[�x9��������g�g��a%�bg�V^��B��V�h�4@�hI�1㙢H=���P��V��v?k�E}����7C�-�_� �fx�=�Z�s��}3O��J/=̑�$����Z�UKH�lŘ�*��__�'p
yf�XF[��2��5(Yf���y�;��aޏ�a^��qs�i��*=!	cE�?��>�!��	9�����j9(.���Σ*���&�"^E(�.G��a���4hN�߁��I�����jVw�cO�1y@!mr� ϿG�*#�Kd��9��]	�nd�>w�,)9v&a�R��c5js�'ٷ>�[�TÞ�6=ӳph��Q���+�̼4��C�_LK�.f�e?IM��^�:m�����p���g���m�j��^�������QYB�Z~�`���li�Lf���$��Χ��g���RU`au	��T�Jc��l�I�'l��G3��c|�jȘjҏ�uO�τ����Т5�SD�W�*�#�cf��k!WF�@?�S�qL�֬��z�H�p5�9_� �P�ƞ-�T�����:�#䐥� �B�X�.X�n4{Q�OKM~Ƽ1i�uԀ�YU����-�p�Z��Oɜ'�U|��ԧ%WF0"�]x�����g�[	��D�	d��$7�	�΄�g��i��֊�1v��z����Z��*�����,���ц��8iV1�WuO���ݛYl�D(�1��ov��W���y�Z��Py���c�m��:�^�B��5_�&�� >���z�gS�C���l�O|�?,��{�Ŷ�bXBt��< z�Ȋylʟ}���\|E3bG	^Iɗ� �/D�{3Xp�۞�8S�B���׋$�����_�P�/@&���B�-J �����>�yj֢���Vm��\*�M�TZ�m��{/��!d<�0�q����X�@s���6DJQM�s>0ف��?����b�������>�����@�Ozm���qhY��$�N���w�l=c�#׉�N���Ӟl2ȗS?�?�?Q����C�Z���V�#����<��~�ㅥ�	��q`�D���TQ��k#s����dI~��=�6q,�%��i@z�>�%}������\AS3��񎬹�2ֳ/m"{���뚀X*��s̅�cP��=���?�d���ZQ����F*S���kc�CF0f��H9�M��Q*���'x�G4;��,�i�w��
�I@��d��"u��Sugk@&�U�|�B��UiȬ�A0[� �\H�|!8:��.�A���C�!#��bȹ��F�U��{�8CE�Y 8�����o��!QS��}O�*X��/^�-$��;��>�u��J���usy»�6��ů�A�cm>"�7��vS�+�Q�ы������ʰz�0�6ڞ�½ #�5�M�;|�u��p+x��ć_ch�H�s��ʡU.�W�j�.�m�Ñ����SFD:��=?Gq��,�u�7A�ݢ=��-V���s)���>TLVϯ�h�_�4fn2���GL�Z������/mj�7�����^�^�.��o���ղ����*�J�̼S��Uf*TgQwF�!��n�������%O��A���ޚP.�����_z̝���~$eY��ϫ��@���6�L��SY��q��n��hG�ՎU��zR���ڎ�<���'/�S�P��$<��S�y�2@7�u���~л�B�;�"�E�=�`q8в͠&�p%Q��ވ+����4U:��H62aNeg2�f�Q/%���#a�i�8����!*�T��g6���b
���22&�s��i�t�Gl�+NR\��Vp�3ܢ�
�^��fx�1VE@f�q@W<(��Uy��P>+�r��|z�d��id��j7P΄�>��Ŧ*���xQB+Ϊ�tV��K&J�gJ�
�ePՈ���,h���(PUyZ�t�"����Ot�V:�%�蕈����;]��]�E�::��ۃ-��h�c��Jׯ�h��%F�IaC.O�R�'N(�(h4�-Z�[i3�v����{��2�]��\�#��*Dk��+󥱫[�y��ᡗoTT빱�p�(�I��qx>��q��ׯшp;���6V"vS'U���ηwU�8�Da������@.t|�V�h��_���H���{�4WA s\%��ǤMɻ}�VP/P��_��
�p�uV�����*�2�����m���O$���t>[�S�h�A\4�-^�}����� ��&��w��' �˱lT	O6�{���S���Q8z�v�G��3NFX��0M�H�E@C�{��K-�y�s�a�WV �J�i�*��
Z��<!��x�/�!��&�e��(=��z�̻,tV��.f"�8��C�]�Ms �'�?��ҬIYQtb3���n/M^�x�M=Q�SZ1�Z��p��!_�5�� HZY�n���[UC�Q� ��_�uB��qED1{�3:�-`pD2p����
���-�x�pv��"ثA��l�{��d�v��	���L>0��F�Ob��������h�Kec��%V��-��">�
qn�B��^`-�A<�d��� �����i���%�8�~ȯ��MK%#�j�:��;��a����r�< ���<�l�U���F۹B���Y-:7?>��x�غD(������Z���>��W��F�)g���'m���V�;�akH*�Dx
�R�s������ag�wa�RʗQ��oC��f7�@��=	���00b*��qܗ�����J���H�1OFA�����f1;a�Δ�	�sR%��I<�Ɯ�3�v-~��t���-M(	�#HNm������V�������(��=[	�*�E�%Sj[3�h?���f��W��}RBY;��o`u �Qt��9O­q:����G�M�Q�������g�&�t�ߟ�-Mɷy�u3�f��u��n�b��V� �|���$$�$��ɢ9�3��%���}��?&+o��|K�6e�4-¼��h�+E�]�7�/Qj�|7�Z��쩟{6j��~Ѓ�B���
��QB����o���^���
�m�.@�꼳��҈�sU��p�|3�E0�Mz2���O�u�9R�q�݂))���/=YD Sf�_L�H~��U��	(���w1����6<1�{��$�P�keZ�݇I��J���`䳞9W{�_��I���mI��ܮ�O���\C���i�Gb�g;�S�ݷ�eeޗ���ĴM�.e�ZH��w�L�0�_+�Nt?JUH댒 �P0a�9���5�&6�E<�#1B^+��Е/�U,S1�ZP���ȣ��&r����/\0;;�ʷF�j�=�����w�W�����DO��w"�sYk��N�(F+τ#���hꆬȢ3E-S�#̖�
��R��y>�43	kUݗ�ጡ���oU^g剞D�ȝ�?G��;�Y/�/���OO���.ܕ��& �>�9w�Ϯ�1���F�TVN�ޠr�cօPT��0����%SW���]!x�TD�x]��jw|�B�_�ׂğ��R�n0,M�b�w�fN�C!�ܩ��M6�(|ˉ�=���������F6&?
�!�cJ�b;�˅�]
��3��Z\�@��1����q��NY!����̐�̝�#�sV���x]%�T�H
N}4���G��4E{�� ���3��Z(:���bY�&��}-g�JJ௒	�n�TLR^��w6��B��L[x��|�a���Y���>�d6�9e�+7��7���_k��vp��=y
~�N�֐�t��!����-ZK����x��LP�A�~W�d�f�5"I��:�BWq4H)",�ȅ���\�L�!��� �[�v����V}X���,���E=�����z✽��m�l%Y�i66\��i��wM9R���˯(�O l�O�\1Ǘ���m����r�K|V_�L���#�e�����I�$�@��u���	d0�R��dC2�+��dvMr�pk`#��O��g����i��x�����ý��J^���|����q����-;~k��%�J����:�Ud;C��T�p�	}Y��NmiL�ޢ�������fɮ�_�%i+�o�$o����bo)�"ƅ���E�@_��_�!3��;�����_S��_O��d�-;o<�W8S�_�}��G!���v�Yf"M�<
�$s~jЪ����AuJ��;��s��ئjA*u>�5�A٦��qg�PW��N��.���7Q*�9��X4����~X�sH����1�".�c$EM��u�����%��.��� r���TU[K�4Z��(��+�g��:ϼ<�5���ˊ�4�����Me����1Xf�"� ���O?3�8�+7N8څ���w�[�S��;���v��xc��/L,
wyS_`��!�M)���-����6��L//�j��Yd3��#9Ƨ�בB�"	cN�"N�^�p��6�:9-�<~_�4���] ��y)��8y�	�D��L ^��	S����M|�|Kk�5HD0���B�&�i�_�	Jޣ��V�&$���a^T1��L��(������E�l'.�~]F��'���t{�υ׼�B .�e���[�K��jʼ��>d�q�T���/�Ⱥ��=��eZc�,"o�`�a
�(�j����;�ZjX���T���q��M`�`i�c������!#�V$C^�Z�B0� ���[�3�Um n��Xy4~�7�漢��>U�#'��0I�� �߬8�H&՜��؀�TL�<�����|�Մ�֞�(�Y��4��;��C�.#� ��Z�X�Va�r����q������3X����P�<�,�@��;2�P��򻪰1�Cڔ��&����;�����;t��TU�,��}��ti��N6 9�.�{ߍ��P`���6-�jਤ��zr �P���ߖ�<�4ɐ�<N7�{��OHm����� ՑkԷ���B�I��C�<��0�g�dpW����r/+*���G�=��FŞR�~j�HZ����)9���`��zr}��,��j�Öwp�V�i9i"}��O����8�j;�.�Q0s��Ɨ�$sTբjC;\*����g�#bT+6s�B��Dޔڤ�����wu�s��^��y8%�(��(���:���!��j$C�>��tN�y���NoY��8A,i�+C)�E�����O��@LױzN��K޴�{@�g�"E�s@砺ӥ Kn���Ń�q-.gL~�����ֈ�����(7%2N�aȕ{�>�C��7�k}��m���)����&�0`��&O�l/?����-E8�����!��&����� h [���UB>=�F�x���`�^!^���
����<R�J�j8���\�E������	��1KFӶY��2� QbDP�I�t~#wD^���;�~���*�����S��$b�W�sr��2O�����D��l�L�Ta�5τ�ю$_2��U��|��Gm��'6\��+�P�-������f]�z|���"ŢНOS:�Ŵ���Y�\����up`0oB:έ��]����U�"ap3��h��j�r�U6����@�pMr��\x�e�4o���zp��(:Anb�m����Ɣ�Ѻ�jj9$�%F�׾*`���;�~M���
%�K���[�]υ~S�s��8l��ۢ�ZA����ٟ����t�iQ�5_3�#F0F����VK'$žXj��ݎ�~(�,u��5+�R��a0�����h��='�N�|eS+�}�8�ۦϗ�v$��(/���Z�i ���x=���LJ+��3u�@?�|}� �l�}Q����x��~.��R�=��"�eە&U�;�b:�&�9#�t���i�� �FG�WtF�a����L�줂�Qi�������ȬV��C�x�Jd�0�[IT˔*ȉ[h\x�j��p�>E/��k#t��@�:�
Y`���۾�x���P���6�L�] ���cGŘ�Z�sbb,�Qi����խ^�|��>tͥZQ�`:�:;��hd+h�]k2���"�=}y����mb��.�,�<5Xd$���!��B����_=K�,Q���_th 9��-�x��?o��]�OA�z=z�j����2�}�B0�y�y�bN�w޻J�Bpꚻ���	��/��a�R&vA��܎_AP�/�,���f����T.��)^S ��3���<���e�'�A��}��n�]jl�b�~�WY{�YR�<B`~�R��E�)d�O�Q��
���N���~����Ɇ�#��U�)�U����o7n]�Ƀ50"�H��=4�d��Mr�%���� �Bw��Lq�ɗ��ˇKl�Y��D��!����8�D�q1{�|ws#�؛��]���OqoH��J	��|b�HS�Ql߀g��mJ���	��͍8 {��t����+T�x�Z�  �boT��
ފp|9���P�{{���Gv���m��� �hW�]-�O�X����D�oɍ��g6}�M��0���>\�H-33_��K6w��(���b����h>����S���xG�2h�T�=�����&�#O銩�Y"k��D�����W{{bǴ#��	D&��2��Q<^�{�l�����	M�����p���A�I�D�6�&B(A�	�{e��Y��G��T�s��
�v|�"=:�]�p����������v��F�&4�=���K{���Z�4LD��[h�z�.�V�F�afG���*���D[���7u�)U5��۪��V>H��4Oֈ(��`��~Q����.�B N�(��5����-j/O�Q`�r14���ˆ�^�p�ᆫ�F=�W�o�0�='u`{ľ�EM�eE��]��
��~@Ě����Dp��1�M�B��!�I��U�8��Xr^*~B��{���k��c�ڱ��(�?��z����R��N�����v@H-�.3�n�-~<�牴S��IkWʬ��+T���C��`iǜ��8�N��Y�s
n�>�3�>U�f�)�E�bޑm!��39��l���f5`�s���|��h�ԞvR�	 D��$����?K�&I�����~S�/����-�sDO!��Ԫ��\�+�,���o֗�{s��Wb��#C����y����������VƌVm�4W��Y-��n�L��d����N:�lz�w�)<�Ӷ/�X;5��O�ɰ*������}�HO{1�Rؓ_�*�l��6r}�����<F�+�,�扚v�s�3TLe�cn�G�`V,�d�C���ϸY^k��8�� �N��xK�	f��Ck��c4Z�0ׂ���j#�T�p�[!=��/ȸ��
5��:R�g����p��R||P�ҽ3�6%:�A��I�����T��5u[}�0��L�Ș�eB�n1G�|�|�-рU���XjPTHc
.Ny�Gz��w�=��hbтʈ��\a=8�. �pz�`~�Or �Q����c@n�+����b�c�Cm�g$yx���ǲ^��]��n�>/�� ��]��!�	?�h�=��6g���r6�s�v, ��|�;��[�у��ؖ5�.(�	&�W����FB��t��W�r/u,���h�[�G6����;�#J�*74����'��[ɠ��:����`����X�,�ه�YP�-:�����LS�����2�_ ~"����q3]�h�Ds�MĨYȚ};��S��L��g��ۡ)�ƥ��/eeN
�} >~����yECV�c�o)�Hb+��|�۩�\	���k:zcL�d|2�螌W�c2�}��Q#踇��oa�#���*�i��AQ�^�w���-�������[K���%xb���}`q!�n�^0�7������=qO��k��^�腃���^j9�$1�96q֫��T36���P�U��!�Tq�[o�����"�������6�-g���_C�j�3����P�_V� @���'y%�s�u4�h��4V���?�G����7H����1���	�� }�F��_PڠL��5�����ag�B�1t����J��X4G�Q���D2JO]�u͡���y5�B��o�^����ӄ�~C��!�ݮ���vx#�g�E�sy�l=D0��[u��Ǥd�ћ���(���`!f"]�OU��
�<��.�w,��xDV�5��ja�J���b~c��&HK}K�����d��P�X��r\��X[�.��� �^x�����غ��CuU�>�m8.U"���3^*K\dK|��Q��8v߉L��g�s�����8�^�+�Ͼ�s.,,t/Nsf�ԇ0��+�T�^�5�f��j3��J��2�m��q���.�T��Y������-�=����&��,jS=
"y�#��Z\Te���� �ش:���T�
'i��9^���0gA���=�ʗ���fg�H��<}�B���@��?�}U�C�u�N������4[%�[4��":P*�*��|w� 繧�ն��V��)wk9��wدj�fъ!ρL94�#=��g�(��S$\���Ӣ�Ϋk9ӆ�1�ai�IMZ1^��B��)v�l�0N0�2VJ��#a�TC庩궈�M�2���v�<s��䇙߮�+m+�Y�G���4k������X\�y%v�7uY���B��N��,�M��^�_Iw�"�a.rX���ѭ=XG��u=9~r�z���13n�N�̆�����(AdB����7�l��P9[C^����c�b�֥I�9���iŽ%��ST�YG�v�ڟ�Q��ѳhurE@�P@�5�*_>��:�0�MKpm��M]8�p�jK���������� ��Yw���] �!5UfcG����"���EsOʩ��~��D�E�������]�~O7�Qc�N�ӗ�Н�%�3!��5;#T�ڨ�Ƌ#��Oc��<��_�,+����*��a�A��t���`��A����;��a��c~!Y	���*�����#��7�^@�t'�\i�@��heH���+���;� hA�#էm_����&�iJ�Ľ�*�ċ�+t�"B��P�� E�ח���tR.}�6;���aN7U�7dYSy�����S�b�Žn�;��5���L�e*7��ߝu��aɲ)㯌4<�q
�q�4o��w�)�&N�H�jx��W�d�;e�3Ƭ⼊	@S��V�3#�K3p���tl8�'��S{��"rl�w"��F ��c����ʢ=���|2A1�Y�kl�F��K�O�T�`��4w�Q�i]fe3�y�Y�6Z5CX�U;:�N�b[��`�#����'�4�y����=$tR_0�`���U���S�z,�2�[�tF8$Ec$�i���@���^��:�3	�bDm��g]����Ko�!�hH�_���K[�)��{5e��Gs�𰙮�����F3����ݱi7ŖF�.)}2]|�h��P�Wo�?6�dc{*RB��0ɂ�l�0�~��#�(�j)����;%9tB�3�kK�P�����s�#��QZ���3� )t��b!�{Z��c�V��uO�`d%@>��V�0b=P$o�j�p�Jh��}�<N�Y�qw �t-㳒QQ�Q�W����9�ie��_;d]�P�܆�r�����,R�YPX�5�;�\͝Du�������R��|np�г��5U�'��
'�K�{��[�#��	�_����8+�C�E��F�����[Q��Gk���N������1��
}��Ivv����"O�n��K;��$Y�Ra|�m�Y�����jr�Zۭ�'���#�Ǧe�r����3���>jD���k2����B0��2���%���(G�v\Wp�����:a�~�T�Q3#�[�S�rm{H��O�'|!��SmBh�3aQk �*����}��O���E�x�{��@9���*�3�|dh���-$�xў��*�<</��nX��Zt!_�h�d���_������ħ�d���� �b��3�e��xe;�9��kq�����蝋e�i↞ެCbH`R��5G~��qb����D�x�g�3���!L��8$��mQ¦��һ�9}��ʯ+?-��NPz��(�Ra���0Г��4�%@c����D��Tr��1S��M��X��G�wA���?=�E��K�$�C?�!9��k���3x���g�O<�$����Qou��}mge��;0vE4!�Y�[�Txm�LDh�Ki���}=7�N�o��X7�����Ft�̈��{� ��x\�ٜ6�wZ &�=����&�eMW�!1~���S���Q,w?�96�|Ug'�0��$&�Ó�H�B	�h���1���޼�ߑ�����^�sh+=��e�Y���������rmxB2����S�ߦ����¬\����v��K��S�W�:�Fttc׶;'.ē��@<9�U���t�+���}��0v���ϕ��Ɂ�$�bAd���yc���%z1�*��egC������9��
^<ܜq���DJ5�cu�mZ�5%li5��C:���ɤ��$�i�M�m�3�6������,;!��i�XL,5�|��j���kT�^vpd�Vr��fp�k\/�#k�r��m��EO�q��ܴ%ym��	�:t\AdO�Q����7�
�k�� O��9U�sFQ_�,F�ݥ?����@ұ$x����#���҈פ��O�o]@5eӏ5�!�#7�#y曱��ĵ��%$�.wl��jz���A��[Z�[{���/fԪ�ՆL�$��]��Q��#�x]8H��Z�:KE�c�~uī�<ׄ��]n8�DV�4�������������h*�j���՜�ϩ�1*Ȧ�$�p�CL�
�(�i-ĕ�G����oo"�VA��Ó�M��!��Z7h���%�(�G�|t��h=pܧ�j���.g����!=�{�`��5���v���f���,���,���aO^�!t&I[Ɨx��Q��f� @^R�Xy�D��}���eS$њ�a�åW�� �vUpSY�_���%�4M��k�����˦���w��*[H��	�h$�~>	Q����7��2[��$�{	el�N�B��Q��=�N��$3���q�|qѣ/I�r�،�hv�$���k�h�V���)8�	� ��S[6i�C���Aa�ȯ���xzkp�|��(�T��SL��F=��'K�ę@<�Ս�XwA��\y�'/d����1��+��8�Ù��Ky��W@��Pe�4���4H&��Ex�n��yW�òD�2�o�1h�b*P1� �Au�۶� �:�����WC����;t���쿐�Ep�N��AЫn�W�HG%��ե�!�~g ���K��xM���^^��V�{���BJ룥z�I�ꩳ3�2\2)i�7�����Ey�bه�s���>O^��`�^露A��Qۣv����k��
A���O![x�J7����{����gLWR���r����=M��L
�kY�Lgm��PW��Iətwmµ�!6��qs��/�����3�%^�ж�d�P�ġ���թ�B�k*��d|�~y,Ꮠ'�S��&�+1����xLd�ɳ�(?ge-���W F��#�Յ2�d�-�Pީz��Z!4�O�Q���J� ^Y�J�t� ��^��Ly���]#[;^_�aq�$��Ki*���Z)���ሳ�Q�v�U�����6�m<��䮅�����J�)���2�{#Ug��KmxQ��D�
Rb�s�r嫧�Q��TJ��?*������Xߵl �2��t_v/3*�h����=�p�kĢe�5��^[WJǢ�C/���Kt�'B�j�؊���+"x" <�*;�ʲ}��9��<qh�{H���z>K(�5�vQ X�lG���Ψ�]�BC�2z�S�E��^Ngզ'~��Ӟ�#�S�\��3Z퓸�[���w0c���Ƙ3޷z���x���]�Y�l�iEi���<U�����K�)���"�a����j�,<�,>�l��դf����{4���h�\Q�	���]�(�W�e�������v3�И���F�H�,O<�-0���l���}�����Ih��!C)�J�N��܆�Of���J�I�F;��V��,
�擭���+�8���be�(�7EM�C|��:P���?"��e����y�f����i)~��䮚y�ۚ�'{��"�6\3���zk��Y��x�ca����ve�]�C91�>�I]�<�r{��Vr�x}�O���2꟦� �IQ�� �#�}��#�_��b�_}��W~'7�77tQA�Iͽ��Ex��r��|k�n�O����HU����.|��Y.O�m�g_=<������8u,Aս��R|����sU�"��ʿ��͓ �Wc�}�[F�7ҳK�0h�ܤ��%�"�2�G8��'�� 4���'���%����(����;���V�x���U{�.ZW�� �_�h�UYϫe��e�K�w����2G���ɺ�=����we�Ǩ��B�&�+ß���?{�
�����gE�l���y6�����5ׯ��Q�U�8d�`��: ����>�$�Ix����˦�:Qv�o�z�ӡ��ܖѤ��W*�A��Yꥄfw��1�3cb.h�2����qJz��RxHڎK ��Z����4^lI��J!K�u�+��YE�{teʑ�W�c������*[RH�n�Jy�,Ln|�N�G�$`|���FO����j0:G�b%�L�+D̋q�t�o�=5��`��E��i%�ՕD���!i�Q΅�"c�'��{�/I���"P��w Q��^���5�n�h�W�x���Nɣ�+Bg��7�5�ˎ�d
����8W����S\v�����>����.�1�@��ⷨ�m���(�2M���߉Z	�1S�_�d�I��p��Z�Z�ܨ7 �w"qh3��j��}A'�v~�|�2�'��8����L}�n��s�s�k����_�����;ٵ��$-Ē��Z��G��CϹ,�f���r���@�TbV,����oR�ݰ)������Y�Q:���
ƶ�?Ѧ{���#��[~����,QL=9xk�x�K���w�3�xʩ�/&H`A�urU|u�0F['1�}����TY����7�P�s'�n����l�ɚ7�����������X�Q���7r~10s�:� 3�{{x:���iB��ܟ�o���>��vmXk�i��njZ]�I�>���v�΀�bޚl'�4|Y����z����iv�����|�?`��B�&��@�]D\�W;@�����r�@�"'p��F�z6Rއ�� ^�!�{F�@��o��sB/�Y��v���������q�AN6�Rs�I�O�ཫ[ԁ�o�!'��=�5>��+���Z0|�<M��7O��@ُ�m��''���'�̈́�6,���P���n���W>2��bP74�2��In刿�%�LH���;���+6:bkǛ+���c���)�#�#�5P �R���b쎶de塗�1jY��^�(���7n��#ݼ���4��Sm�"��N/�"���%oP�\�FO?A����%�F%��1�����i�5×��A��"OK"�M��i�p�&���D�������l�Y���yh6%�͎Nj'���s�\�C���n�\�l������hy��߆�! ��5�t�]1�/��k�-Q�0*�UOp���������6H�h5�)IG��UwB�Sbz��������e�ֱ�j�t�;�W�Ȑ������	ԇ����d|�I
��K)��t3���t��CoK[�ѯv�~��ͫ �j��Ѷ5���#�~�������)��x��`� Z�E79B�����2H�40�э��`�^�~ݖp���W	�9�S2�� e�&Jb��-�O��k�- ��h�d��&��,�;ED����4:�~��0;���R T	<�;w�pjl��4��P?o�^=!M��o�	Կ(�����2dJ�-��}v���5�X9}����z1��H�2�� ^7*���]�u5�V/{�=�t��4�.����ʙ�\@u�S���!�H�bzϤ�:@H���M��C�6^I��LSM�)��rv�����|7�)3�*�7v��1��6*H �{��i��XQ]SX��^��؁1naQ����{��P�YӸl�a�W��]���������C^�@Q�t:!�����=B:�f�5��256���ph�;6_��ʥ��reZ!�m��0H�Ӝ�bTv��6�?�Vp�	�8����Y�P��n
�����ص�َ�^&���E@���4�V�ٜ��7W��zM��%���<���G�oLAI�"v��S��tf��S�q��u.N�0��Y�D	S��c}��@�r ��k�N���Icz�Ð�
L��i�@C>sQ�����y���������	�.X��;�T��&��!|wXnJ��^υ����Zd��M����"���B`����Ur��H{'�υ�&������y��~���a��O�0��#J⻎�nƊ�8��1��+����锳[�s�r�U'= Ig��(yaR���l±��w��:$�-��V|�M��e�t,�ݳ/����M׺g��gXw�TL��:Z�K�߆���6��j:��>*�P�r�m�^fZEaR)��ظ�Rݎ�պ��;W�}m��/칝��d]�GUP��վ��0�^�~���Z����e0��h���hhA$ ! ͞�.���&�M}[�f�-�R��ؠ�E�c�Z�TmY_��\��I�f�D�����W����y`AUt�n��`�"��m�Kez]}u�r�۝�
"�a+����v|
m���͕kN�p�HM�Qp"��`��:��,%�M܌�[����/8i�6�!4y1sdz;8���'F�cQ�N.^8˻�3�/l&��cD�<J�c��$ށâѭSޏ�]?f�#o?��C�"�����ʌ(��(}}j��LդT�s[�,o\ą�ԋsv��S|��*Xݥ�Of2��D a��J4.�N��`�*4�O��8X����!2��e��(����d�ex@��T݁g�I@�ҹ��4��`�V�RYd�ԋ�xDp4��b�aw#yi�J���^M���H��N��ꚛ� �9TB�ٳ(W��id��w�$|��h4��q���wL�4�:���AFw����͎��d� �-��T���#J,T�E��}2Įsǽ������K�n(߽�Q�v"q+L�f�ƶ�vu1L�4�96R��)p���}X�&����R"��;���LT�u����o#��C%�Ł���j[)8�����|�d�矉PT�9����+��^�x�sQ"�b�;�����[]]��>�k���s�i�#�S;B���q��/��H�s�k`:<*� Oէ77�ˎ�M�l�A��Jω�-�خ퀧�DгC��"�#Lu���S��ޔ��x���������\�%�������9>�I໤,#�R�D>���1�ծe��Du���$�<-��͍��VU}M��LaI����y6�Y��'���TRV4.Ғ�a���&���R31>eX�����QV���,����;nC���ڄ@�;�%�70L�f��i$�'�jVc7a�x-�)�7����h�	�� (���u�C�l��~z0k�_DE�)�J����nN[u�o}������w
#ԈֈO�)^����a|@ۡVz�C����?oKυYF� �\jOa��U?ߛ󵥗yL�l2_q���߮������,��}�����2M��:R~�J{���I�96��% �7*NJhZ	�o�<g�X��(�<w�6��FȿqB���d��AKU^؁��\2��-����U&6Y^Q�h<����!t*����.��>�am�{HܦDrD��]1�{����'�/�[��=z��r�:�:�Ԕ��W���s(ROC�&(��eU�}LO���r9v�['��p�{O#V��O6?�a-��Zg��n�!rD�y`o��-��]�Ĩ�� -u�4N���`2�ɂ�%E%�(2U��g�H^v��DZd޴F8
�?mn�ܽǍ)��h���e~�=��Q��[�I�N<�A������m����w[t̫�T�xH��	��Pʫ��φ�b�(��Ya��=�I�jg�mw����ih�(���#��_"n��A�l``Y�и����w��|�@��8124���eb�s����������V�M���x�4�aI�ͫwB� (�d,>"�W�WaȻÁ>*�����a�u�(�>F�e��ا�돟�L-qz���{nj]�[�:@���d
�NC4���y�f���3"R����Unn�I�u���A!S�\�[.dS3�O�h��2����e�`X�A<)����n�?�F�-�K�4*�j(�̐y�h7�$@�Fk'�w�MIlɪ�Ej��@:����6ݜ�KHE�����or,�b��4��r6.�">Ѕ6�ժ��=���A�^K���K�UE}��G�R�}Vj|��Ԩ��7]D���X/�U=��)��^��|��l�ܾ|"�ᡌ�^3�%�r���}�G����8�/��S`�t]����T����q9�W���1-�T���%!g>k`H�8X�i"��?ej�8�R'���|3��B�C�u�{`*x$Ax'�KF/g@oA�vָ���"�%"�ː�[����{�3,u��G|���p#�'�~�&W����q��n����H����ȉ�Itk�e�KS��b�e]QՂ�)�L��[�Ʉ6� Y�L��*��-�����6�}I
cu99�!ii���+�^���y$J���HK� F$q���F�k�t���3�ҹ�@�{��"w��/EgoW�DX�nl�)T��(T���j���>�Hk���F�F{�dU����÷Z�20�-2s֗!�Z?
_��׃y�o���A.�ҽn���f���{�u���+w�8�y=J���_|��	�,NdN
�Ա̧9*��E���9sr!r)x�~��R�\kPl�';��qP�T[(�>#m�4�%\]�Ϡ ��N[j���!gq��6�mk��؈&
�ё#�j}:}$�����҈7f�5�<{e����!���Z��7�羂3ԣWm�_�v�\�Z�b.j(��N�>�T���Z��[�@�Lo��G�f'[ä��*�n+W�U���L��+��|%��Ʋ�|��	�Q%-������m�dJ��P��erA/�Z�c^S����c���e^�a��į5�W��~���Kc!��I-�mT���ǛG��a�E!��Y�%�pZ�tgJ$C $��W9�i,�fd��J��6���:O��^ʁ��u�|5-(cF�_�F���b�j���ez
G�*!��2Cq���)z�W�ɻ�a�]X��q��x����b�!. ��%�l{����r��52ȇU�� 7!#�ƾ�&+}���:�Qah��J��TFn��đ#���5�Z���؂��;�	�1��}d�
CJ���Z?����p�/[�M���tVXz�k�{[ћ����@���ºz>���h�rm��~�ofq���,�P���o��R�|x���'=��pw�qӹ�mƠ5�0ܸSlu����W��L��_��C(�MC��2;	�6E1�B���O��V���^\
�m���'w�?*�69�!ha��K�\Y�|A�^>7��C"M�yH��G�&[�Lqɵ	�3?p��Hn�D�!���Ku�{6|`�,�&U�SfJ*��FZLS2�
[^p�
������ݨ���>�ѯ|*��l�}����B��M�x�j�T�w^��gVr���fk��,�w��!r���ܹ����P�^H�u����F�`�#�Qj?4S%&m�(FL�����
T�-gH�����i!
X�\�b���X����->֙���.�? �OcEZs�������>��LF�I��
x��Ԙ�=�l2$<��P�y��� �/��_1���ѱ����-3�45ey�S҃�iW���ա�\�r�ǵ���P�2�D*Lqg���jc�H[E���,�ȺJ�Ry�Φ�xEt�^��d��WN�G6�8�Ԩ�0p�Ԩ2��b�Q9������^�/��uoslX�e���(5�*�a,�z 	\�J��T�:�~̽X���Xª�)��9Gy���2�"AP����/v��l��B��.3`j8/�H���vDIwF�e��}��[�z�F��]
�� �W-��s@�?&1�#����P3�OA�`p��P�:Yܧ����\g��Ɗ���v��=lb��q��4l�b�mL���(\	L��W�!�H/�I�1v��F��v��z�y�_ּ'�L=��=+a/K*q�0�ƙr��ҌH� :%��$ ��K����鼝x���P=<})����Lk8�v��pN?�2�ǌਡ�%6mb?f��Z�����NZ�B����i��MU�Pm�4�9Ki��(��>�h�iJ����a���u�'�9Y�#c��e�MF��D˃x6�/-��;���K<��9�oh���5�
[b�g��
�1�ڜͱӌX]�<雫?���)m��2�\<���d1C[�#l�/�è�۴�/��5�W
�VC�Ր��i�q�DNm�c'�̬	H@f�(2ڣ/���T%�h7BנQ��t}�t�+��]V�e>fz҂�t�Q�	�1jj��
D��}X��%��MP �P[tꮒ>[����W�}@�qJZ�l%����S9*��Z�b␩6���q�w�FI"�$v���|#�Z�S��?Ge/N���XYQ�����E��AF��	Q�����{�0���:`����~z~��m��k����	._�r�
�Q��q���hw�%N���!�#�-C�o����&�� �O�"�b�;{޷)�Q�*z@Tȧ����4x/-�N[�{Ǜ8��m�K*Q�fO{����W�
lj~, q�hJ��.Zy��\��ѯ~��ݟ��;�J��r�pۂߙ���3��E��0wIV���gɫn�<7��I��ʐ������;p�U�{þ����=�R@�'��iʇ�W̃3��Ě	mn��?<vߡ���[����+�j�u����������1����@?�g�`��QA1�U��W��v���ĭm���I'��� �FuZE�xtk���z2e��"R��>����2�k���V���K���~L���B0bI��욨:�O���ȿ��f 7j�:/�����<,�#��ؽy�6o�ύ��q6�7����,bf��<g|>�&O�����۾\�
��P�v����,(ڽrh�W)��2O��sjk���@��]����#�;Lº���9�otR�W�(ri]G����W=(�$���wTؓ܅���W�S�T6Ϻ1�p�Q��t�^�`t^�Ф�뇡�~�0�<�e�����*:��1)>o`�S�5/?\a"B��5���5inȩ�}�E�Nn<|Ci:Umg�j`�%�/� TF~g���V5��W�c����3Z��:^q$Ok��G�(Sٱ��F=�٬��[������G�T��ޫ���>,��p�,"F48�{�k�7КZ�N���m����x��?���V�훼|����h�dvh��d��y��a'u8����Y�����F\A�!�	�o<���4h�pF�\q�������ځV�-�ߕ�n����h�J����;�i/�AX{����v΅�}�P����DQۖ��D�^�{��d"�Rb�i1�|x�M˂����"j�u��;��"��U\����4�y���^�c��|_�#���l~�֠Y-�S�������d�XKH�	G�/��02�lZ�{�g"s���0�7���^��{)�o_�a����2�4|��D6�mO�8��pU��ڹ��A��B�� ��+��*���'�ߝ�������]5}�/
SG$E�k]22�7QI���%@�d���o�h�.�5;䎗xr&���?kH�p�b���e7GyC8�,��i��X�"]��F��4���X4���y6Pz�� �fC�}��n)�:�v7�������n��/���\���w$���&�3/�Nx	����T} �N��c/ڔ�k�,�!�"�C_`/c��h��arMJ�f���Y(�ύ_X4�g/S�e0x����2��oݢ�+'N�k�9�7a0nZߠ)����>���.��j�^��Jf}`Pb���c�e���]q�PI���0f�k+�����ף�_<=����1�P�@���?ػ��!�Q�_?��m���N�NEV )����z���4�� �;��tG���%���N�����GAU�T�:T=M�Ԇ�������J�EIz$w�F�F������ ���:�����~��5���R����x���m�C�������t���oG7n�A�-A��D�M� &vr�,2FM��%8��Ѡ������H((���vf����8��c��� ��D���~�J��/�%���ȷ-�l�т9@U�%���|K1�:����As�5��O!�qO�zb8�d��ժ�勝��+�7�P��XE0lWF��'����?�����B5�g�%�@�n�^���/R?���G%��+���	��z��N.5��� 	�G��45�P4�z�߹��o�ʭ�!)�Ǝ&=Uu;8s���y��X�ϋ�jݺ瑪G6���y�s-�o�f�fE��ﾴj��*t�ʱ�#��N�ei��G7RK8��m\�o��n7��E�����=���t�k��H����ow4�d�,�Cc�J)}�a,�X��'�41���A.Uσ��ы���E�Vå9;zX�>�F�Zk��k��n�ɦ�8h�i9��������B��L� �@�(�V��q����^@l��*ʅwtt7��RL�t�����]o�#s�̈́.,�F�M���{jQ�4C�\� ,Hj`a�vi�1�-�q����
M �5񰜵}WD���$���SqV|t�5�+x�g,Y+�rF��Մ뷆n@^�O_���V�6g�^�0�mkC��p�>f�Q�Oj�M�]����w�O��{="&3A\�����m���d�	-�ͽ|<��X����E�>UD��(�v��!�_�Ff�-����c��0�|�˯����񴷝�����7����E �֟qR�縯6���Ϛ����`�6N�2�7.
�QH��H/��DJx��S<��&�0���5���*��Cj?B<�F5%�PB���]ܛ����y�r���G���Ġ5������*'�*�_b:C�c)%k��I����� �3�{�k7Ѝ���4��� >��r��~�6㮍JR�G~J� q�Yy@���xa0lu��=�Ch��2�Ka��=E������'��@�>�0��?d.�@_`Ng�j�Ub?kЖc�����m��ї��&$X�'t�����u�������,�$�%�r| �
E�&�*�W�BqQ|��\	��ۚ���!@mXҾ쫎���8d�iS�u61Q��EɃ�6��0~�0�h1V�Ak��PrN�4��J(�.��X&�ړ{�i�ݺ	s \#�G��l��+�GY4�f)�&ΰ��N����q�ƻu�B/[b�BB��%�m�:߶kr?��/���UQÇ�g�gw�������S��|�᪆N�AV�'�������r�h�Ǯ�o�����E�pH�_�I����pr64�!��S�ts�I��VEJ�S�x���c � ���K�����*��,(��o��{Q���!n��ĂF�XNX��Ǹ?�����,��]{)�"�e��ߟ���$/����)<�1�RNL�P2l���)�!���n�s�8CG� !bHյ_�r���U��c�	EI�u�`�����orB^��f��Y]��=-�P�7�aXv���q*�|:@@���%�Ӱ5\�G�@ci/��d�b;�xC��#��&K�o�(��V�j_܇V�RʸH�Kɕr�r��~�yAg\8�y�v���J��^��O��Ɗ�+]|M#1�8I�eQQ�.�q�l�Lx�t�QY�!,�K<����=�N��m1gT�����`g�M�j�F�b�� ���b��g�|WT#�� �p�{b����H����(�{�����-9�W���>ӌ����1U�-oh���xAibcG�-ܫ�!��I��i�v^8�*��9i��
w.a�Oq��fx��V=g��XH'�˦�����V<��#�7`�ݓZ0��U}�>��}�*���o��]��Vo�`��F��U�i6�/�0c��A��O�P,��S_>wx�ޮӡ�
9�ف�t��b���+Gvމs'���^�Y2d��52�
w�1�
|\6��C2��6���`<�{��1k��kܞ��,5zy�������Q���#��6s�ŝf8.�郡��4)7�g�1�i�ۗ���٫���9�=�؝ �^�����>U�����ڍ��t��~�#��j_E�.s��/�<�O����.�gh�T��6�%��	'���2M�����Xb��".�kn��k��d��5&W��z>x"Pȗ�*�Q��D����tތzz�-�;"%`K�	Yq�������@'Vb��V�א��^?e�oЛ|b��o#K2���s�1��/S�uR��K�na(�<
g\��r
�T�p*�\�ǯf�\�1��a�n�~^�G��3n����9;Yy����B����8�aPvFx�h��o�v�
 !}��\���A�&�V� C����U�'"��s�2{�<?L�F������5��0}P��hqQ�#����4'�CA�&�e�~47��\Wf�c
���r��)��e:PGE��Z�][�Uv�P�D1.������NqY_�9%����HÉwӢ,��1���PB3����纵(�1q�Z��*c�������?1f�c�!�O�oTŤ���V/�B�Ʉ2�m����
s�]�͈ś�o���cw���y�ȳ�H��01q��,�G ]�]�2˿����ݯ��*J9׃���%F對��۟���0�b��R��S�n��|��{�@{���
X��0����~����]kZџ6���U��D�Z5�(�š�"G�`�/ATF�� V���=(�o�P�ȋ�n��F��+��wǞjZE!�9^g����T�������ײCŭ��N�Q��A8DÍ��k�pǮd�����袼��G�T��������,H\^ ��A�`͝XU[�E^�҄[�$ 	E���y4���A��7�§҇,�^�����B7X�&�UGJg�ۙ�V	4�zC�pd6i���_�ۺG�0(E+����H��c����1���gI�8,ّo�(5��$7��a��Ğr�;��ƾ3��aU��6Xk� ���J]�������H��`ڼ0Hp`��I�y�ie/ćN�����É<B�����\����]�.��*Ji��~��Iρ�9���d������ڹtVs�3������G����M����ꓷ ����ҡ̅8I��0���
��;E��3Q���., !�z#����,l���P;)��o �H�T-���1p��Y�&�L@k�(�<NĠ��`�Ye�B�*'����ݤ�yf�AE)��D�?r���	���љ��o�$�|3���p���O"W�":;�,;W� ��:�0'��$�w47�y)��uz@T@ J(-�;����w�%6p��5&�mn�Xv\Ł�
}n���%��Du��i�Z6O�4r�P���]`��HI{8[�Ju�<���H���5�&�/���am뾈A!�F.���H#bWd��B/�w?XI���5=ԃ${�'
�`\�0P�*�r������)�!���	B?L���1���~�,Ue��=dA�7�O6�ԃʩ2c��%���+��v��e�c�C��W�F��͢�_*�X%=T����e���)��L���!I�.�g���� ���)�fa�&a ho�n�
����0Tc�fT��X��x���q�D�`c+u����> ɨ
!A(��{��9�/E�DL�V�nr�!�W�Њ���Q�*���"i-^s�BˤH�����<�J����e�[�Z���CtHi�xnatQH�R<8�a�+�"�w]��@"��	}����UuBo�-��J�T굏g�ye(�T��#DT��.��?_���!ktU���TLsl�:������rat�H�PE,�Ci@h�g8;��Y8��(#���jz���|W*X�	$�̥D�i+����j?��o��2�c���B����1���}��*r��5F��nT����<"O7]M,3*W)��>p���3��y�l ���2d�蠖���&%�dK�6�ܨ=)�lQ�uh��,��/L��'�ʆ�fe:�7\��4t�hw7��9��vQ��g�o-q��D�>�������.�)�:�;�e<	`��5�~^i�O}o��tH	#�:/�d�)�(L?�a&8S`���Cs�ꢑ�HK<�G\��g��fCc1֯$T��2�q��
�|牳@8��Q1juӿ���V��:�g�����b��%S�Ұ��l.x�Ap#> =]�ۯ2�z��
��Yg�s�D
�[z�5��%}u�5���d}��b�K8C�Y�Wډ����_6����`����#U�!�5�n�硊�0-Nl�k+���(�mF��Af{�a�{�F��3�� �n��:$a7V�9�~!�U�.��BC⾃�?�}pV�Cls@�Z���%� ��(��]��x^��al����>�t ���B�9��'kq��Fj�;!u�C�yA��:v*L'����),Xu/�z��,�O��'�d��!��y9��x5g�kw��%?���(g.Ǣ�8z��>�2�@��g��W��)%���7_;Ģ䃊�U����\ZscI��w&
b�R�O�εHk��?�^��AN�'0�#&Ѻ�Z�{���u5��a7�fX�gO�C�lq�Y"
xa���9�:���[�jwVyl2�\")�����`��~{ᙁ�%P�w"\����[���^H/��h�`[�]~3:���;���9���N����'��/���աAA*�C"i��5��ήhR����W3�>+���PE�
���)]�	�����
��	H����J΅!j�6Z;QF���{��ִ����	q���V)J��g����ةH��#	J��ó�u�F~����}F���7���ovZf��!g[�(����n�gWwp1mÒ#5�5��G������
~FV�x���oȒ3k!d"�tSl�c�SW�)Y�vٓ���<�dT]�v�HQ�V9I��zEN.�F ��4�o�+׹-=���(�$���>�>������7�����nf�,)4�B"��l�ݱ����\9[�w)��}}��:��jΕ1�u������4�lFݵ<�?��SsƓ��Z_`B\,�ڛɢ�]�.��R���&<�=��"��]����<����Jy�r"�����G;]#P;u����©V�{��ͭJ�2��BH˓C�4.�S���]��MǷ��u�IMl����S�&{4�懶yȘfH�?1�_7�duK;>ڠ!�mHp����o1�S=B^r���N��5������v�Q3 ^C8��T�(i-������@Qu3����ɓ`��32I�#S���3�Z.͕8t����Q�5x2�Lrhj��	\#�Em��<83�yK;��[�޽���B)�g��,=C*���d̥S�k�Kvf0��;�\i����E^$p�1�V>Y��%��sͳ{�e�|��O>z�~p:��p���?Q��w����惓�kkH������4ld��p���πe��� ��V�ʈ����he�#��8 b%��,�5�R��m[���H+��>�;����e�M�G����ǦD�>Q�_'Fj9��BU'��A9�*�ݼ�^;��H�'�%Dr)J�+"��h�B����_���;�8^���� ��G=�(��g�M�qr!O�,�܄B5��Q����`��c�6�H�qa�v@Z;��~4hJb?�^r��aP��f��'~����=c�d�c��NEB�L�Pw3���K���N��T���#��X�Բ�^!Fɤ�VyD����� jEa�F��5�GڢqUpd@}q�]a�2���4����a��_� �=��C\�݅�6���@w�5����(9(#�R��7�QR�SQ��'�3FwI�v<�S>\���W'���5��urR�m���B��Y�H���ͣ��`p�  ����Uf�p��m��vX�lɩ �u�zZ�+&�R��P�m?���xy��N�{5��m�B��z9C��./~�[E|� n�vuђ*�{j�@V���b�w?�t���Q#���4)e,�VI�~��N���'x���&!��␯%-��Y���,���� H~)�N2�<������e���KB�c�xդ}/W8�6G�#/Y�ԙ��J"6+��/��[���#���#�?�����fyN�������g�?l�x�,C��[�C}�\��є������Ǫ�� �E?Q�ܞ�\T�`�4��/�)Y��/�+�����v���F��I�Lko[�ȸ4E/hB&_��7x��J�����\���  �둚I1���=ѻ��)ZgŊo�ٴ�T�:H���� i���t��SɎz��r穇pӥ�f�mL�a�[�e�q2J�XG�n����x���O9jƙF��YW@��֊�؄8%�L�4�����w&��
~�m�G,t�JO��	ȿa�̻�*�3m�e��Ig��s�)�m���h4hr����߁�~Í$*��n�����l-{mT󒦥+�����m�;cEc�\�����>괘���}�o���p'�S��d�p�$���5N?ɜO�i\��e�f��L[y<��K��P'6�eK����\m3���s#�yP��@:>�e�$�[�G�Ӻ��S����3�&n�ӝ֌���ݔ�D�w��R�BVlQh�����+hb�Ao-L+_��F��B�c�o\	�>E%���lP,��t/r�]���<��I��Z,q�
��F�_���ue~x"�7����`_���-8�.&��q00�Vy�j��t��	:1�\�X^[J�����rU!��`,�>�����(�ALQ)Ѥ�x�2�X��&���X��+U/`RJ#�[�n����.�u<�B�t�$���JT�J\A ��Y�줩E�-���n���A�
�B?i����>�7��6�p��x)�D�#"e���РEԝ��W)}���S�T���*kŌ��/W}0��)M#�1o�'����h䋡������V�ҹ���&�0+�]����ϷG3t������ ���a��ˢ�C{�����-+�`)�����z��~��S�n\��-N)m�er`�lpQ�J�k����g����ɵ�.1�R�=f��L^w/��;�v0h��[&p�v�4m?}�� M"�'u����]�5Qޒ�g{)����aoD�k���t�����)����r%T��F��ǚ2~�����aRK�����b�!����w^H��^����v���̒+v����� �rpX�<<��8��A�Ϭ��c�q��S`� 0�Эs�L�ۯ$o*R�K�6*°��t����F˩,#��o�9<�*�.I�e��@�
��𴨰s��6��T�O'x�"�	���`�
��Mԅi=�L�k�b��셣A��Xuԏ��Ӭ�<�KG�"*�*�TG���5��٤+��>4j��"]nh�a�N�8��BS�IT(q�WHA���*Qv�:��,����h��8�C�q�v����!tSǘD!l�jrqZ���@�*`�E�~��x;��7E�ΰ�6��$��{I��^d�	b=	��/��ו2Ź��%�O�H��E~%�3Ȕ��y��IE�՞��ݑ��r8���
� j�cڑw�+XJ�%�1�M�Ήi�Y����g$��'C�[���`D�k�f=@�F#X.lKܹ��2t��j��^w�o��٨��0�^�C�g�Ɠ�~B�QA1G��������Q���t+�L2#:�����v�A��-�<d�1ٞ��7�mK ��q4��\��gN(dF� >�ne�"E�>~���rT8� �)<�!��"��K-��������l]����e����M'L��4y�A���T=`���z�߷�9��;bz��j���׼k}��_O���|���P��E��ᝂ��'��?�7����e��l�f�M^������R��0��\�w1���R������u!��n�z���5:@ 54�V�5ά�FYz��p��Rcm�%h9�<��B0�_c2��/o�2�,$�'9��=�.�,�JS[݀C�qV��*"i�2��S�����P�]��^���W^Gܯ(3#�@�ݣ˘0����BI�5��ĊK8)���f��v%�o�Tc�ϳ�T%W�
-�6�uk��~����ŏq��\�3���𹗛I��l[�� g�
�T�܁H�
ؒ���5l�g°Y�q�.�b���
���S|ބAS�0e/q1��]�&Ei���B�V�����6�X��Ͼ4��X�h�ON��02�c.$F�1�^�����P����˟��� .'@���Ou�۔�բ���Ӵ�f΋���bd��/�VV�ҷll�A�'��G)��J����G3τ��1�pQ���ǖ���c���L�2b�(�n~i�z]�;#yk��
�IXxت���!�*?���[Ly��=�)9�A��w1`��H�����cN�m���[�`�܉!@h�
ڍ)]�G)���T��z���`���IN�[{Jd!Da�JMs�w�ʔdgfy��5��q�46�'a�M���H��F2��3D 3�,7�=��GD����
�i��𞎭�Ae��G/�R5s�pO��;p^�%�e��F���r��0@�G�u#/�GB���N;ے.έ��n���0h�c�� >�A��.�ʂK��/�j��v�S��L�@'?��x�-ǜ�~�|���H��9�f��5c��G���Dc+��}���"v���~Ol�b���SF�0���m�aD�����+��$�p�J�[�u�����	�'�+^�Ջ�X;Ϊ��]����������8X��M"sɊ�9K���'D*�D�b��"�Z>�A1�2�üM{����D���'\y��8�7�_�>t�]ϗ����@DQ���{.�H�"j�0F����ܣ�W��'t⬝���	�֏�w[����fB�M��I��`�h��'$^	�mu!
*���n� ���A7v����{�֍By�]�Recd`�t���������7>��@K�1���zJ�FFQ��ث��l.-�T!T'����PSN�ܡpɌI� :�~�CЉ
I�+Z/����޶��ܚ���~��5:"1�����3���>;|T�8���%�M���D)u�%ūM?�g\iuM�*�Y������	n�5�P��k�}��	��=[�R�k1��̕�N�'*���Ms�N�Ƞp N�|@�#\l2.�u�p~� <lu�v�ȗf$:d�?9b �����
�r�1�|#5˿J
e꥟�=_�$a%��gK����h=�02�sÛ:�r@H��5�b��ܓ� ��ZT@7�V��m��<؂�۸hL��Ҵ���vɳ�M_p�uhE����ċTX�$�0We�Ő�2�2���+���&B���p&~L�X���
|�c���r�;-�Hc�� ���͆����8G3s�U�]i�5�UdA�D_��MD!���C�	�$���%��e�x������P��9�t1Y?�C!]�A.���n���V �w-���뼿�n�;jh~�Mb���bR��b�r��h/�ٶ�N(&D��9��W	�p��顥��ݝ�>u��`[�:AN�'��),_�Mz������O���a��bU��,Q[c�����f����X$N�;�)Gˮ��"�Pb/���O�9~>�U�;ֶ�&ӺϽ�-+6I���l֎|y����_͡m$M&�a�F���C9�0ɛxU/�c�"x�i��^'�v�h���e���z��ƭ���Q�qC1���ڞ����_��~V6D{U)��Diq���a�� Jr5��ɟ�b6�2���:���.��[#���Kj �eKh�����~c`�8�sD��52(��w��&�P�gԧRT���qP#/�S��L��7�-���`ly���8j�W���C^&�8Ȑ
ey�r�a"�LY>/e��~���]5���:@�e�&�1�`�/,�"9���u���nސ�[=�o� 'g5��$�kЙ��i�����h߄1P�2�J��41�š�7M�]�US'�xSkX�� 8&�=�~�������)M�83Ђ���X�0++}�cW���V�^r�Rȶ��,{-�E"Y�����'�3
T�o|�s^7�;����}=D�_��֪+��'}�fJ/�TC.��no<d(� yy�q���¤z�w 5��X�Tq'Kʅo�����d���������Ϛ�O���uF>����]X�����{p�����K��:zJߛ��n��+q��02.�bB���T��JK �q�֕<����Њ�\|a �>᤾b�g���DYӎż�sw��}�n�Y��d�\��%�1�����~�M��sz>P����4��A\��Ţ�+7q�3����<�
�(�Dޢo�\'�j(����~�3�����.�G9�+�Q��q���TҤ��WILk�j�n��4�ܵ旨BO��u�a�y��]=}��랴�u����j������.�`�+N��}��``;,��fh�+zFB��~%��5b���@��_�:���>��]�}��s���h#� a|U%�^�����V�l���g�p���8QQ$!� #�r�����*��[� +Q��J[���d��`���tN�#��}��������S��>A��o��;ha�D-@�--��W���;>�n{�w6a��N7����!H�U5a�����u5������I�>>9�Ї���`���,��ΆԘ�}ϵ\����~7�,~A$n�<�̺��ы����A]2��1��v�w(�hyDɇ��S�Q���ς�WB'���i<��g�	��X�F��m��T#��|!$��?���t��}s��Yy���xo�{0�gB�d'�aR�س�#fQ_����H�@b����ڒЯs�p7�(��uШΆ�)|a�c��G���,�sÀ�p�ʪ�8FCw���K�c���9�����:/�eo���E�=q�Z����ϑv�e!�Q�&�ua�;@�8�^ұU� �Z��W���C���$�r��؊H�>�:�G}g�=[��#@3�/g���xN�����9a�Ǭ�[������R���k=˟��q���0H	o��>�[�3>���0,��+Z�T[́ģ�6<���j�R�ꩳ4v�`��j�~�.*@	P�t�[7����?(��r�[�Z�����32�sR=���%Ѡ���-\.��#ϿPL|�z��cU�e�-���Z�8h�s�oFY��y��'���8�S#�b?ӂ㥵ϔ7	�'<f:Cd���ҩ�V!�q�����Q`���|sq�".��B����t����S|M8��6r���`5���)���S�{�3Yb��%<��9OCʟ�agE�{>d3�%�h���׉c�:ҝ�����-	�l�O�|7*�[|��sJ�wگf1��,cVĎ!���d�~,�����{���j���@�Di�-��A(2����0[��_��������ǫ�Vi�.4搎g�V��"R�#���n��N�'�g��h��*]�7�n�C e���v1�ˬ�����Lo6�d���Z���ȭ|�(�h*.��SV�[5,���)��x�,�Ʈ@�O��7��X��y9Q��μ1�����R�Ф��?r3hm���dOj��u�E{����tQh
$��΢Ѹ+͢A뀭�8ß{N��J���0��:8ps0&���]צ�FL�g�;jMk)px�x?/	���-���ij�~=�⛭k�t�.�Q��:�g\���v��W�f;w͕z�_��hE�6�?�*��%�j�����B�YT26Q�	�+�����ab|`_�"�D���I�X%�b��sm8�=�bvs(���O���7a8��o��Z`^�j��A3zO�GM^+Ƣfu⚽C]�l~d�ZS4�޻��y���	�/�)$#�ù��s�6����tX]��O�6��9�E2���挻sY�V9Ό���5��,ˏ�����I�Ui�(j��?�b~$q�����B[��re� ڂ����0B_�]D��d��
��;�J9�[�>�����
�������gؼ�\S<�����E#�w�Iҁ��.=ZmZ��w@(-��$�e�a��"g�0��%�x&aG�^�N����T] UUn�2D} ��ˊXH'�!�k�rM�pB�����~��e�CB��� �Wg�B>k$I�7@s��U��҂F�~��Y)����m)ILR<CˇcN-CEԳ�G� ���BԢr���9\�__�bߌCGc"���˂�]\�X��RO��U�����n�(��
`} ����A����t;Ĭ�����+h�H��`�=��c�=Z_^`u������E�N2z�m���ň�gxߝ�w����bF��S�VO��^�'���b�l]m���sCr�C����y'�[٪Z#M��VfC>��!&KK��6��n\��E���#��J���.<P�@������	KɔP��7tF�8�ojG'4D��~�R"�r�e�{�';_�ϝ�*4�!�C��'��-{b�.�_�d�j��r��N�Lt��Q�A�ά�=��h������d�nř<��:r�C{�W���slIl�}�t���t�$�0�i�ɯ鯶�6ҷ"EOS��l�[]��зc�s�4(�(p�h�7a�#�J�q�Q�D��w�e�H+�bJ�� ��m�vx����Ҳ0�GJ��>����n2����`�򵇷>Z�ˤ��}xV��=;�g��Y�ıs�G�UZ�ު��?u,�ƓB<
X�#��D�����j7a�Ή�r��4�G	�!`�e�e˜w��܊�eg��?ЅX�拵�%.X��H�MP��D��|}=p���Q��
x����&Щ
(Zr(�|���~֤��J�Z3mЌ����a�_�����ʓcEk3���"W+��p�������3i�ݐ��Á�tU=�󎩵�FQ�5d�sp@M���?�O��|��b�qt*i�knY8�U�ȑ���~�\u	�y*�w���k%Z�I��J��߁Rd�Z������x��y�r��e�`23�"��t?�K����f���O�W�,3�M"4�I�>J�� q���������U���V ��b�G1��c .��k��|+�ad��f��{�����ЮsR�Kqܔ�)�ʂ8p�
�4w^�A+��#��|\0l�GK�a/����tGt��Dq�9ޱ;	���/���ro
�7��e�ȝd�[��G��9��qO��s%����H�w~�Z	��żNqK��Ƅ���::��^QL�} �B�>�{���"[����*,�m���C�o�劜�hE�80��K��)Z�ڗ�Dv���kHz�c���*�;����u�����m��ܧ��Az����:ۢ���k��`}:�~⫍)���'����E��*�5��ƽ�q�w���y~���ys�堦�z�/����N��yTE�g��)��yO;������p��<��ѽH��*46�ٓ��h`���g'Z:�DYr����wT��T:������o>�ٍ?kIؘ5^4��!~�.4K�|L� G�O4Ŧ^�,I�<��^����(��r$U A�+<C7���e�V�K�7Z����o��)>�nV� ������,_�g�p�3�t܎�uV`��SgL
����u.��+S���:�m�f����
Gܰ �#+F�֙T!n�aq��;�J��YA V�@�?�4I@��1N��H�su�X������JԢ�7̪t�m[���E�)F�(�+^Kޯ�X̏�*��0�L3�o��0W�y�U�D���u���"��A�僱��t��v��4���!�g~���d�A9��/%},����J��o���X&�6a����"U����������H9  �Û�H�:5�3���7�AkL��7��w���+��`1��f���kDt��p�q�61���T�u[�����\�(����kGr�[B�YAG�$%�<�y-���q�5���i�ƘHd��j'�x�[�3�̦����1��!�YX4���hN�G))o�a�WUwg����֠�&V�MQ��˔b|�$w��FB����Q����)�j��">[�{@�ukcG5�x�6Y_�*וg;�V���4�T[�)Y�����5��hP�01XF���]��vG,lJ���R�D�����pݥ(����WN��.=`���n�����qAu��A(>DP+ƧyP�p��T�s��u�V��B�j�h����V���d�!T���T�)M���Aע[�a�K������q#|�G�X��Ơ\'%�S���`O�"q�ɰ�1�D��8��ա��._������sZ���j����r"Kߝ�xq$�v��O���`�~w����/nk��!I�g/�`�,������ֲ��0QZ'�"��"�[�gy��* ��5�0���;��0�F]'�Ti��X�2��
��+*��Jp�1'�m|lA:�z�ޔ}�B��g�e4.)y.i��ށ���G,�@����K�.j�&S\�� d��ΛW��0�85�:��bJ �tO������{@\��'b^HV6�4�(E�ۣ��vӨ�y��V��"�Ģ���d�شX���	����w�z�v��zѦ�'��'��m	�|��S�%�i�-]Lqu�"U�jC�Uz��lbh2��ö�K��f���{b΅�@)l ��0x >��C��n�5�����u�Nj�5�Z�T7B���;��㤲��ʲuF��)V��̀WN����q�N� k�RF��S�vf��c�\Wq�&��$'�(�y�1�w��P��k����2�)���B[��Զ�d|*���U=����G�v!�<ݢ�vN�Ї�7>�e��D�	�0���t&�ˏ
�˽!��~�!�Bo='K,�z�	�4Gmo�z?;����Q�h��0����f5i��9PF���~*}<�wD�W�d����Lsˋ�/pOu�)mt����]��;L�����6��3!HL�]�Y� Q����2YS�rg�}��`?7t������Sa!�g��^1n��_=�q��5uN�Ҝַ|٢�!S��n�qA���;���j@�a��T	gb���z�$Yo�jQ������_�ha�0��R5���s��:T�J�Ї��.��P��	�^����J�`s���[�QRBt59	Mp_V{L��=ocE+%��܉Q�{]>���l����U�p�a0Ǔ�n�J�0s�ap�'��A1t��v>Y��7d�h�טK��:�_�b��DZ�6NU~��}>���\m�(_��S)W릑��L���v:Rd�n�K����I����e�ɧ$9��9	}:�ԙ(�_gB�Dء��> �a^�8s���"��2�o�>�Rԁ�f�"Р"+���ݢ��}�w^<-�	U9Ŗ��-5�:�{F[0��٦����y7gmr�w�X�,�/�;��A���܉\<�V.Ir���������ef<M?�o�>aHKH�>V��H���W�R+���(�O��x��QH�d�+?,k��)�&a9�;��ˑ�J��]*�e�f��$�s�p>��W!L�sB6�r��^�<�"kQ���	�_X ���<���e��Z�w���X��4�����Ӟq��H�᪺z�U� �hرFF�aA��"����Z:E�Ƃ%�[D��:��.���E�g40�N90���q'�Dl��S�x��8�������@�K	�E��幗�=j�S)�Sx��n Lv+.��뾙f4^I*�-�܌�Q���h'A,U�:.�cWN+"[�#�kІ:� 3eF�Kj5^k6���S�%z����(�L�z��h�!|�~e��<e�S~x�.���s#�6�I�d��ѥ5����;����N煢 �F1S,~�!�W+?ٺ��вѶP��"��X���dW�6�Zi�Ҧ��}l7��*����qf,~f݊(����#�M�)�|��
%A�aխ�Yl4*�j�/�a���^�/�������)��}L��W={���s'[.~{-�@�Ӹ���/?�׷w��0{�O�F��[�JF���ՓVuq�z���S"h^�pM�'ЇH�Eq��?-KvYB��A�J��_�G��$������<�Μ[�ڨs�?]v$����ֱ^:q7No-��'A⋹� �Tx�Dp���Ĳ\q��.Dn�6�5,����UJ�̍wDL=���ŝΒ4��k`��O�R�}�Jq֑|�`�"=�����?@�4N��e/@�Y�q��E�FB�;5=�>�_Qs\r|*]�eN�P�ߡ5�1��Sd�2�-W��~��aܩCX#d
1+�`Gڒ:��g�z��y;U�8�����7��A�큒�9�QT�� I�eR+�$Y�oa$�y�Q���_�jnE��lee���B�WJ��W�=�m9�{�+p������jv!ݐ\Ne��Z ��1����4A�Tm�"���Df����p�^�Rt��ǃ]6ɲU�s4�����I(af�%�l!@Pݛm��Mp?���5����[|_[�Lg���o]����ai�.W�>p+���i��-|�����3��r6�/w�l�y�&�k��b�S��uv�B��hn�Bs`�4M�Pk��R+"�@/%�{�����2ʪ
�a<k�{m��Ə�:���8�S�B������ad���b�G+۹)?�	���{�k�#�k���U��C���8`�קg��V�7��~�X��uC�&2�+·��˲��Ų8⺡�pn�Tg��n�^ڨ��N����H�+�̒L��~@|�㞰y�#�2�옽��=��;�߶�Ɖ�*�7��ɍ����h?y�ZB2�]X�{�a���&�ŏ�T8�@fm!�fI.A/�2����s�� x��Z�c�\�Q��3	>�j��c%���Up�daJ���W����]ݴf_^��K��[R�?^0�;/_����/�X�uǀ��j5�h�z*��cR�τ˧��a�Y��������>|7n.����E��+<ó����SI��u*BƵۂ#��F�{�Ԧ��M	r����P��-�'��2ԃ��l[��]�*���=���0ڳ\�-Ehؤ�j���6�s���j҆PRy�T�}&�����l�垝9���&�4JD�<]�u?P!��{��*��ٚ�J���q�����Ͷ.D��B<������w��jy/�r�6���,u�CrO�M�A«�����G��@�1�wl���H�if�hc��΄ �"h!�Z��+�y�]��h�jF�����:R����<K�n��JM�~��OFuY�$aK=�p1���wU�C?*���u��J['4i�d:�s�zSf�l3ve\�yt@�,�BB�"[쐑�cpC2�g(3^���g7�Q�v-�J%���5�x�<q��鐱Ĕ��╖���_=�T�?�G�l���4��,N�[y�G��T���ubw�"e&s��V�U��ݲ֦���		I/T������~(��ז�w�������m��Q����1
'.�Mn�&������n��0�,
���~ަ��G�3B������֙�6�4�i��vk;���3k�{�Y�uy
��������=�ؘ�1G���h�Y��s$t�9�	�-���JQ�$K(�bP�!2Z$�N�r7��ӹ������qS�BS�ă�����>���@�K}��H צP����c��V��S�Ƒc���p�ڶ�j`��+��f���U��l!G�br8�#?��7-g!�mH�1�.�R� ����6=X�ï�#�@�v�f�IvU���5	��Z~ƒ"D$�H�V�_�݈w�Ie� ���YD��w����uX�#�� ����G2�����^5%*���� u�?�M8�S8��Hk�7������4��闁�@�9V��1�Wq��'b�R4e9���S/�iv�˶G�S�-5�fC�!�M���K��T�ꫴBP�g�+R0����5^��hDW��R��.*huT͝"���G��ta����c�6��=%$���U�Z��.b2�SA�KyC�����
MT�M �N��%�~C�e�+>�b�2q�l�c���������A�\>�����R���G�Jc*��Xt���H��6� W�]�[�5ƥS�$��Bt�M�ã�P��B�w��FO�Ʌ��VyƅpY%�D��T�˟���g��[��'�I�����%��@�F_���P�z�8�Z�tq,�t��QO����_����}�+s�)��3읔�O�dIJ<;1^TjX\�'��6���FzL�:S"쥹���d�ִ��"�'��	:$NӋp�qy�R��@�ؿ��?�+��'^?9�-K�`�{����)� G6����cs.(��1b[����ڻt� Ƙ�f]�L"a�d�4���?B���'��}w�s@�rAk"ь��Р��~��[�ە��-��]��ѷ��ӑ�Cu�V�����+�S�|Qq!�����.�����8?j��0;ϛ���;)e�&�`�WgƟ��,<N��*���m$r�No!{��Z�X��l�'�C���Pc�/� l��"?��$]]!(xh�T��
*�p>���f�=y��1�H�����K����c!����%��N�ȑtq�&�׿���>����KN�r��\�|��:�#�=i̅)�C1
h�56��)�O��\����J�谁͞��A;ܭUl�Z��%����`Hؐ��_d<5-ê:�W
�Z�r�e
Ѩ��Q��\��F�Ś׺g�%�����_���R���mB�����X6����߫liq!2�b�@�Ԍ�'�Ua+�G��*�X;$NW����	�,`l�]��U��V�?����/�Yѳ̯�'`ge���ZiYn�J�r��Ev�ԵB�3���U�=��-�����|6����lU��;*w[`��ۉ\`�����I�(�S�3k���sK�'B�ܫl8�*$���ϰ�<���H.��:�m��3v3Kv��D�*�?��}���o'������-��^��@�P;X��@kL��-��F<T�}��RSt����ti�o���eqkѥ��Ţ���&�v��	[\���E�R�-�����i�^���w��-e�β �����ֆ��+I��_P���DfUʊ�U���24�0Т?�C���B�:��#tC�ZN���˙�}%Z��2��Ze�ŋ�����1v���)ɴ��*>�\_�vy�v%�4x�k��N�ֶ�HB�`�-r�±.���D�g�Jz�j���8a�n��ת�O����%i�D�damL��D�g��6;��@ퟍ���� SsXiG#ɿ�
��k���꣛���Q���"��嬓���s�Q��cM&�d���e��;�7���P�����ɬ	�	�G�X�����@�H���A��ן�{b�SC�i�E��m��3�E>)Ep�8����������B�s4;[�LZ1�u7��)b�~3`.
[�C��Bڌ�GU�f����U�i����g�����4p�K�'�^�P*�-��u7K��պ��,��>��� f�lZ�*%^:�[%2��6i�}j��ɒW��K�)���,��r��G�/���[p~^��̬�BM\��!�Ap{�v֬�2���'b���w(X�륩�t��[m�
����>������ן��q{�e^اdC.�3�M�L�a��,�H��P0F��f�q�l�}��oKM���&D�� 9ݬE
B�9���:K�����A�v<3PU��.�SҊr�a#L���w�drZ���OiftWE�*�]P�*�&C�>���r�~~V�ީm��ܿ�q�B=OA��?�'�e�*���rC�7��}�A���N-3��l�\��G���c�y
��;vԚN~�Μp���n�3�&�}/V2@q3���tYJ�!�A�R��B�dn�a݅9��y�z+#@)���3�y�/��#o�(H��
"���Q#+��ˮ�J�wD��c���S�h�8���n��ڻ�}+N |#uW�OL�*�{��A�ʺ�||�˿�}~&h7�߲���B�_b��9a���r�*&���LOnc<�W!a��s#�}y��%��$��[B�H�:��F�['2ʒz٠@u���:�.d�^���f���D����x2u��Q6#�I��N�����_�c�$c!��},���"�v��f�"�-���HAɫmI��};�Y��*ytu,?z�����)E��N���7���Τi5�����qWb�o2 kA�W�f5׵��r�A� t����q�qHM��'~љ�Yc�ެD&�~� �~�pqB��+E�詀`��{������F�0k�$S�M?�Z���͎��}6��Q����;@ @(	��f}���
m*�`�Z�q�������^n	q>t�[���H��a"�d�'��щ
׈Ų��9����?U69$�4�+肌��H�V��`�9͏څ������Q�)�80K�z���b#��Ás�|[}޽U�����Ep�����3<e�n�cQ{��J�MIb���Z�L����&h��]و���h��_,���lHU|5���,g�^�M~�t��ϯ�C.��j2��I��b� �Xl��k��̠`�xJ�E�����J�}��
`6�Z@O'Q,��"')[�P�1���Y������ꞎ��	�S'��,=v:I8^]d��]��~�.(v��E��K7�9���g=`4�y�HG��*]�m��:H�����œ2_��\��e�gao��F�,D��,2J60s|��h4l���<q/P��`XX��-VP�N�6I>4+Ǘ(��G�z�3��O0;2����\�;�a�MsҶ�=瞁�+J�Vr�Z�Hҭ�	�+��fk>�p��B ��ǈrc��:H#R�Ιk�,J+�d�`Ɵ�ݘ(��T#�u�S�������ʟt\e�6�P�O#��^T]_ھE���@��G�r� }n�e����׊�1�(��+�h
t4��<21��%�ՊT�.f[�
V`��b45��*���6�(�җ�������q{X��==RD��ǥ}��X�޹�!��V)���"����g}Nqĉ�a��9^=��a�3�_�q���m���yQ�n��*M��@%h��G���E7cȦl��Dz�cl�Z+Hޙ<ؽ��+.�<��8�ۡr�M�����+�y���Q��msIrK*�]�$�*)�W��;"��ȼT�Nf³��\����gm����3�J�D�ϐ�a|�_��=#n1��q��w�'��]I�fq��I�?�|��� մ���`�E���A�+>Ʉ���7�5\����-���G��z�_�K�=O�0��c�1�L�L@�~�qd�_
�x_�`�4�x�Fޱ��_G�cH�W�ҡ�O֌��g}}��h��� P��ٷC#�bW{���11��2\��8�	�=���]�Ռp#9�a�1�c��e��~7%�����~t(�[�M��R���í#�T�&�����hA�����"=�ݪ�2�2���H�񷃟��O-�q�q�/�c�)��Őc�k�27�v)����"܌���{�������q��+�S�F�l+f�-�<ȱR�"�X�Z�i2����0�r4�5�N�Ͼ���N��&Ȭ���(�㓯�x%�����G��0�5�ɸ�.'T	��_�vPsσv'�jnB*�����O�*pH�-���p���Я![)֠�t2���8�uӅz�|"������{x�%�`͓]�>�!j���U|�x�g�U��%lE�2
{�q�oz8�am�/��`��yD�a'��7��me�2�| q
���	��N�ê�rH*��0A��B_�B���%����J�D�E�:9��F|���������hC�) 
�6��(x'������(�@鶧�}���Ǳ���ޫ�C��V��
�r�����ek��L�vt?��Nm.#� ��Eo��lSc����աUn��h5�G8�������m��j+�<��sYoi�t��*1%
yT&e�!��
\"�y�� ��?������dԕ���R⎧��dH��E�P����G���1�pE<^�ڏ�'Z����]��:����3(*zw9�y���5]=������^�eMM2RB#����t�BqQ�����S_�+�K��H��Yl�.����e�?&gUs贫P:F~2[��W�"��K]9�C$�*b�o.�N�pV�M4�52YC�HrS���i_��ͣ�o}�J�A�Ц�\���� �SU8ph#�����7��]��*�B`�9�h��Q*�{s�a=��F�໪6e����6cT�0S������؅��So�1��Q8�k�L����E���X��I��̕�M��oݖ��R	�	���j�ų�Q�X����{{<���p��|��#�b�qQe���E	������;ih�{M��L���(�Da)5ul�=z��� �4h�}�=����&]5���p�^�K=��ʟm4��1�yiOO6m��n��9	�k��6�9�QX��h�q	t���/��8��]�K5�Hc�n��
�!7^l^��@�P]�$Y�ԉ�2�x℉���hT! ��ʌ�����2ʗ�D9O������j�7�hA�&�ק���=_��| �E��"L'΋�:zgo�ɸs�R�0L�-S����S�	]ԝX�J�{�N<f���>GՀV�e�w���1Ί�4�YXA(��, OF'���I<0�; �̆��$ ��V��@|ҩ�)����%����|)�����򳪇A9=�_�]�A��飌g늕��JFi��Ԑ�Z�q����)Z����X�sZ_���oSed��~�g<��~�
]�������<�q`���d+&�);��5@�P/[�X�f;��5�j�����]J�OdUs�v�|m�!�)��م?j.8Fm������G��x_�4p���M��Q;H����K.�$"���}���
�ʾ�jC��EqE[��F�7n.ZV6mBv�$p�~�ܡ�����2����%�����$e8}�Q#R�#f��F�~��KMם�	�z+�ZS��/W�>�}��f�Fh�7��]O�4�힙:�X^�����xh���)z�J��,����]{mAyU��	Q��p����.����}�.�e�9ߕ!Ù�"G�>vF+&���YJ����g*K���(TE��+T6���j�w/���p �o���-f�N�,6au�^��_�7�NS"8�6}��P=M��t���߾�����s?��O���^"|K�(��We�ax�h?`-��r�� �s�v�.����@�a[�˧�o'C�1�@}}�W܅ԖMJt/�XX~��۩<���%�1$�ߝ�;c-`�9�|���z�
�!����o��;��b`)�q��^�ϡs9]=e�^��*%���BhH��覼�@Pq�A��D6�uXvE��ؗ���}�1����RY�\tn��6	;�Qs����&ܱ��ډ��)�����O���KP�y\n�^;����������$��P�J81����|Q��t���c棨����[.��~�lY�@�G�����Ӆ�A�^.�|��`/�ݜ�ޱ� ��7���#�s�t�S��r*���*ؔ����ɗQ��p>��M� ��#�M.�M%Zl"P؝[�o(k݃�3� ��#���a-v��^�5�/T�Ah3��(�4�˙Tڗ
o2���ż�#�p�~U�!���0?y���I�Tsm��0e-��^�z�s2����@��8���L����ڌx6���8����\VP����d'���OD�&��/GV�W��ҨF���PB� ���'���;�:���^�xk^Pl��Wۗ�X�1f�	LXu����Z_`F�~�>Y�K���P%Q�G�@C�=iv�d� m,�'�<FN�~�(D5�$��9�Q�L3`�Ot )�āTd|�Z�_ �J�x8Uݟ�~��t�Ԯ�v����d���;�IJ�T� ��|`tk�#��͹8���&��g�d�wz�� �A�2Ko��"v�U�
cJl�(��LIs��dN�T�Bb7��ޟ]@�ݑ�?�������g��������E�V��F��?ݓ7�;9To���&ÛP���龊��!i6�"͚���9�7�T��1�`%�*64�Rd�E]��Y��2K���Jۃ�8vx�*����* _�q���$��a������,ʦ��skЀ���l7����v�FS5M�����h�e%�]i�%��T�H�T����BՏN��"���2I5�5�}K� NK1�s��Z=^
⌌����cD.����	k_��2a�W�ҲW��m�1���.�I6_� ��$�˨��Q]zv"������|��R�iD�Oz樀.>8)ߺ�����T��M���VF�z���칃�Y�#A*�x,�ւ�2 �x+�Ö���	����[��ᥭ֑v���G�r�>���@p�y\sOC;����x/��,WfS�?�y�[�K��	y�� .��޻��28� ws�oT��<�R��/)�� �*�����3��.���H��V�0��O�{t�'eg_���� v�����ƃ�u���Ү2�>y� <�>��t��kMq(u���P'���j�I+D��`�ӳ�*�d)� �9C.F�x���=,B4�&�������)�5l�5(c���՘��ț���R��u�U��A�a}+�p�����ڐ,��_�ƚ` K�L�I���p�{�Ќ�<�{8��[_5��@��[IR+�Ti����c�6,�_�*E�b6�?jVm3����x"ͺ�4L�pvŧ"�F(3���p���� �?��<r��6��i!�*D`z���:+0�|�+���@�s �j��"������C�H��G�K�'�8���̼d���p�^��Y�)�'�ί�	��2�N��?"�%i����G�D�H��
����ޝ���j��#�	u2,�ٵ�1�b
9%p���V��j��&����4 	d4>F�CӦ��k���v�x跆�G�k�L1�I�=}꠮��Dg ��p���0�hN-؉q�8�3���Nԙ���6~�̉�������6w$�i�����f���n �`geB����[�-5fs������w����v = ��,��Z��Im/� �������3�&��l携sQ�,�A	I]���d���T7D�%����qj�ɖ�P���vXZ���#���1?/EUװ�QW �H9��W/��/��
���i��3c�E�E��l���25�^�p����P��si~�e�'[��Ǎ��ԧw�^���k7IF��U�J�_p��T�|�$�J�xUAFD"=׻q2Ka��W�F�\"�D+���i�IgS�k�B�ٱ�r��NN�of"{'��^+� "8����~������!�}&�p��y9�9:��!��Ur('��;9x����Gx�J�V��7�W�o"�G�G&���#$�[2��VF�xc�d������p`+���8�L��y��2�~	�'MP��c^v�|��L��0?t��n{��ɏ����V��%I�%%n܆hF��y�����n_1����Sa���c$Pu��=�J�n�MW�\�+k;u��T����<5��7V$~~9V�a&<�qR �"|ƥ��dZm����'�x�<�Qiwe�7�Zt^1�P�O���Ms����69Z1^E9�>}�B��vyJ�y꿛�Xq��2�|�}��2(0l_4�a�Ҝ���67䚱Qޡ +
����ࣗ�l�y+�e��ԫ^:�M�5_9,�\;I�[mnR��B)��-���~֬oL�k��ǉkΊF�b+(\�D�]�êT�zW��d�Qux�EL���nT
��
-@���r�2�ym�ӳ�W���R��)܀aS���	����b��L`����pg���ց�� �����Z4�p����v��Ʉ��G?m� ��7D
�y�ШoNWһqN+�EDzԟj���9
@��X�\A�%�[	�������*�����`�jm(��|0�V�v�����|����k;g�WX�o_��'�=��?V��X���MA�n���E��8���/�2�+5���n�?�J�(�Ǥ"i�եO3�DkTb��� �x^ �v|�}���(�}%5�H��8����X���}J����J�ƭ)��iֽ�C��,1�<[�>�>��	�>�K[={������G�τ���W�� X��gm��5k�`v�^n���5Cg�}X�awԏ#�� i������4cB�hQ�?t7PZN!��Oﾘ�td2�BB�����!�:�)��'(���A+�k1c��z�s
�n�5�
�# N�w�!��΋m q]��1$����q�s)"<�mM�wY�7��w4����d�b=KR�v�FsX�fI�kד�`��	_21�(�h@d�}��i�D���!$��tW�yq4C&�o����e�F��x�7J�ښ��C�Tc��nd���K�\]���`�5�s� �_��@�sޗYW��$��O*�ȵAO��e����p5��q���ܘnd�$�� FlE#��l������36���6&;g�k
1֤����&_Hi��	�0�駵r4��Q��2���j�����.�n�~���w�yE,��P�D�-*�μ�E�g�l�}��U-���H�ta�y�f	'�c�XW0cV�%r��~�U:��	���)*����S0j�*���ZmP=򆋩V_k���C�z�U�N�p�Z��~��'	��^ؿ�~2�`lm��Ý�������p}CB�,���3U�QKZx�1CJv�R�\jYn<��mb�j*��w��9>��}�?�K��ఈ	9�&�tx����m��B��4����l7s��@�n����OR�@5��((rd8EM�6@X���(kd�&_[��Ǘ[�>�uZX�"<
�m'�Ն�D��7^��7�J]����w��(r	��`��4�^��ȸ+�pS����2+����[�%h�]{L���y�o�ۅ�G���R�v2�_D@M+� i� ��c�_u���1�jq�I�fH�_ec�L��i�X��D�hwJ'mF״��<(�]ĬK�:ŉ���v�j)k�i�"-L�-6�k�����̭-W�ya��ـ@I�O��Mʜzub�r�w�r��ɫ�.��9 V��f� �B�����,p�:#�a%Bjg=�ӷD���;6՘g��	%y�^<�:�m����!H�7)8-H�=ՙ V��,F�XQ�c5IoX�����ȧ��Jh���2;J�⯓�\�f'Ka�Jg�R�BSo ,\?����n��:6Z���h��>����A�y.�Ћh�i�y�c6���M�R)���~�4��'�D�w�ywT�ϭJ��
��(j�2�C-u���
U,���)���N�`z�䙚6��/�(#��cs�y�'�2��i4��W#S~o(h��4Ӄl�N�bi/�
��6�ˠ�.zQ����:7'<W&�s]_�)yLi�e�	Z��$sRs��S�,Qc(<d����/�
j����lVU�ݙ��?9$�C4���Rr��A>�fR�Ůd؛���3�7����
K<�"��ʅS4�/]�J>dF��t{��(���Z�_�o��`�D�Qu�AZ��yK%?l� �\�2x1�F$�����M�*(Nx����4�|Lo��u�
�|��yI�K�Q��~�
75�G�e`�R��[��9�M
��3H����ue�<�İ�Ι�����.hp�`��ݭ{B/�S�W7RA��d��x[��+g�~6�g�~O�DB���ڜ4��_�V���*�$^�UQ��N�c?ɥa�����w6�P=Yρ���Sv��s)��Z	��Nf�U0��;r�{�H�e�?�6�pQM4,z��&�$R�F���{�o�Z�Թ�H0�뺧�X��[},����6��L:��$_���^[C���d�!��k>�R�� �~6B��Y�Ej�b�;�4(9`��nݜ�}�e�ڕ]>O�ЫNAL��hE�Z�H
(��?�4T��
���.�PZ�}o.Z�p@xb	�p��m��c���E��ͱ���h�a-
<�ۭmJ�z��!E�U�G.5�:�y�tұI��X��D�E���l"ol�����Q�}��X(�[���l�c\�U���
�a@_�Nó���� ��/dQ�ߙ�e�Z(�෯��K����Q;1�t�L�d�F
)i��y�V킲�Y�%��� ��˽���t�{U�($؆��+��p��ƭ�6:�"�s\r��`��_��>vHb7�%[ud���C��&9��T�Z������6�`�~y}����T���!�H��qj���4$���Ԥ^R�ٍ4��2J��M��[;t_d��2��>�y�8��	��7P��6��&ϓ��p�� �@s3��DU�}���������Wh��i�������u�H�OG��]�r�5+�~SW�]pF��e��E_Xb���.�0������1as��R�꒝^i�#O���]&/ 1����X;4�=V�Y��"I3�Y���|ƿ[�3>��!'B��=)C�;d�� l۶<�,i��`�%��"�}�2m���xx׽��V�|���p�1�WB�����q��7�m�Z�b�qzy���e�%V���l��ٌ����7p���U~��$J3�Ry?�¼�����NRS*��[�����-]��,�J�팵�zy֫�cx��r��9H_����7����X�9a�"E$iv`�`��;�����]!ұQ�=[�����7��U�rJ���*%�^U��$(':�v��C\@ƅ��u�"�fU����f���plg]��B.��h���y��ψ:�I�V���I	�N�ݦ&p�<�8��b���xZ�E���ZU/S�_Vb����\���D�>0I,�(���LaU��H���`�ԭ4��낑z����W�:��딸��G�Ϗ�Hl�L�����\.><B��$	*�K�<7�e�3$�1�9����,�^��G<�ؓ�7������'mS���O���כN$R�� �i�z(>��7+G�O��9>�A)�@��.-�d<�t�˿��R�\��f@0�x/�/�l��S%q'^���j����+c��>P�O'��GZ4P�M�f���R�2u�]���r|�>0�Ӝ1h0�Q��ns����`��[+.�翠T��yQ{ځ��`��l������;��>�ũ�*d��Q���mh��1�hPAZn��P�&+p?Ey�]>Y�/�{��+�!�ڼ����%��u�Z9���V_��gTnmo���YX{�n�.a7� �)E�E�?[[�3��w�]��َ����׽QB'�\���°f�%���9���4�m���V��P����뙹��s�'��"�g-�O*�q��9���m`���k�+���?{���],'SLX��v���C�W��z0�|4��f�'�-�iN���S�0#��9v�N�CY[Uխ����?���W��ݮ
 %_	{�xaW�#V)_�O�D����\({�WƲ�Nh D�6���hr\���e 	�7IU.�l���C��oa?�*���M�j�)��l�*�spsq q��dݢ����8��UՇ�G��xŬ���=K��$c�zt�}-g_釜�^)9�E�hg�[����������X��ӡi�@��e~�l�6u�
}��DT��546��M�y���{~�I�Q��/p{M%9mn�/������&�R�[b_�Fޭ�U
-�sd�_��n��y�A@��Ys�Y[���q�R��2���nJ��Z��^o�{mD��M5� ��~3|��(?�����@����&��rW���CBf��vv;U�d���Eb�B�;ٙF�Sv*w[�{&���o�����%���p��=4*�=L�\������9��aq>׀����2e�ԃ��q� �����~N='(�X]����cPd�nD�Vw��q���B2�R�!kۍY#Q��7C��_���mb������[�D
-��ee]
c\�����V��q0�,ـ�l�@޺���r<�ź�}\%���|U$=�x��#b$�vڸlZ6{:����޽[�Y ��͛����[O�ҥ��F��oc��ෟDp!���֞�n]�X�s�B�����e�>q�6��]��p�M�E@ZF��>yFO�EVaX�ܵ�i��|�#��s���W|}� �(�I	@��لB߳��L����*
��(�s�Zf?�L�=k0�#�gI|���}E!�o��[dJJ�DXf�&�T��<e+��Y�q����Rkp1�w].��AV:��m�Ôcv��7�f
���x�D�V�9�B��0�N	��&e�{�s߾M����,:_ß�����4cK�)��d�HH��k1�`<��T�^~�y1V����������`U��dEԴ�ep���G�T��>(�ns�U���TB�E��-���v��.��#�Q�PA�hZ�Ss?�[�Yvm�8~���ӝŕ6�����)$��)���s8c��Y�� ���X���'ǘ�m/��(�K/���mP���"د�C)�i?��U��ج��hI�5�֣�߸�U���3���²6F�j�`a�RC��gz��Ҹ4�H�\9����c�8������!ο�
 ��5�e�J��=S���?HL�Ӱ_�b�%g��tl�"0>IR��/�6SZ�硉�b:�'N��ZJ�lSE������@�X����\��{-|�G:{N��UΝ��`��`Q(A�>�"��@7Lm08�a�U�K�:W���8�1���I&+�sL��ǵ14�m0�p�;M�|9���Gax�/*�.�4u_o�����%"��#��ke#��R1$�I�\�4����[x9<ů�ϔ�2n ��Y��>=�OO���L,�s ��mtDb,Zlӆ*;�X���.�yͼ�$y
��<'ydD�*r����)�N`�V���k�H�j[�T6��%��{�׌Xɮd��Z������k����Sl⚕,��.7§/����ܓOn�\t�Il�̮j�8aC��ROF��M+6r��;�p��|�w��2)�[��˙g��V��}D_��9hZ���Տh��/���j�f0c@���1{]�T��� �,Ei�昽Ct�䤥�ny�l��Xd.��xΨx{��}����*�qq��4֠1����N q���?��#���{w��Ml�׳��iA�U�u�6�\2�)箳;�B�O�����S�1 K��1�j���j��
_�>5m�SM#A��Ѧ�$u)�[�} 6|�XT����x��|��g�Y�j�e����]c�O6�)ۇϚG��74����XN�P�%��Y�CV�8���$�v�+�	�S�gn��gp�O������g��T�Ww$�;U3l��iB�͂gT�R���E�+Uպ>�����R-y��?Гp��U�!R��?U�SY�|;��c�?x��8v�](���:f�ss2�w�@w�X4�j1�Q��-2v9l�PDQ�7�'=��S�(��&!|N�
|;�s��[���N�V��r7daFXq~���KSm��D�UznY�X=�L3
�F/kn��G+�H< ���8��k��Kx�ݨ��MeJG����Ӽ3rI=��@�X`��� �����kj����&���\% tN��q�5/]���M�N�{�AP��Ƨ_ L"�
��`_۰�M�l�h׭#������G��N|l@��N�Oq�BK~[{�˘�u "���΋���� �>���F�B�.�q��ܓ��m�������*`�tO�R�����J��z�2zؿf�~��;`3��z��~Nh�?L����]eD @��6&'�c�u���&cͼp���q�D#rU���&@"l�RM���K�� ����-�#P�B��r;U��:	�,8J����2�J�H^��m�#�PUX���_X7�҆|��rU*��3?�w��oQ��H�7�C�����/1[z����7.=3�Pa{ҏ����<�G�ޝd�פ"����!��<�\�,�?��4Q��t|,����ty#�L�K��Yp�.�5���;�;��K�,�8��F�#��{�z^�N�>�/��z|��^��d����)]ҳmׂ���I�S}z&nj>��rxl�?�<ѻ�|�Á-@���޸N�d|������m]�$x��- �d�E	�B�=�/ ���w�l&6'����F���sy'Q��t2{m�h�O?� ����V���S���r4r6K��-��i�پ��/�ë�o
�9y<~��e�q�H�re���w��LA�'8 �\[���-�-Xn�m-XlYy�������͘���h~��n>�Ϩ+�Py��L�h��|�9G=�	��`p����@��u���C$����&��Z��:dvl/��s��7�~8��,�h:|�NJ	�n�G��y�Eʜz��jm[
�-	*�����Ʌ��w0�Y6	H|ny�������`��ܕ�uVhK�s F�����3�-j4t�G#e���{���'Y���������6���S�y;��{⼧kw�Z�(��ч�:�_�}è�fP�˥�^��O���?Vh5���Dz8���ϥ�م���ms�!��[��ku�L}.�x+����:�Ђ�OA�)D�$��L$���÷=���]����Y{~.p��<T����ˬ���Nޅ�,/�� O��n~��/�KƳ0��x�k`�������Mn��m#!�a#���m��	Rǐ�̎sh�d��BL4�Q}y �lq��~��j���r㗦�l @F��,���@��dR�g���m�VvM����@�q
��̀��?���=��A,V}|#m��`p�{Z��Hu|�~7��������wX��5$����4��D��R��>�é�͍�#vࣉ+`YgՎV��j�	ʌ4fy�W��h�B���v
�Hh�Ak���(,��O{qn,�!|v�l���~�sٹtY;������x�O�8U�w`	/�����B)��*\�~�˻�钾b�l�R���@��{ge[�3�.�0��W�de{�G|���#����Dp��Dm���|�<�,$�๸�̸sJ��ݸ�#
��OO.��0Wv��xzҤ�L*9�#�61(���Є������f��� �/hS
������G=�oH������}R�ƣ���J���Z�(�j"���?����q�R��s��\Q�/�6t������m/�j,P��9��P����t`uH�G�4�$��{n/M�owp��M=#J^&�l-W�v�,�����.;C�Y�)�.�8��}e��2���?v�(2bP�'��� UUa��i=s-6�^@�ߏ�).ĺ+�AHi{c�i���ߋ5�r�l�ֳg�I�+^�QF���Q��9��ܝ��K�x;�f�9P�0>}�\�5^����	mn���qjM���ܗ��\I�"�>�j}UJ�A����� �N�|֎Qh�aE� 3�'�-N��]}S�Q$W�|�k����v�D�S��փ�/�$a�]�d`����"!�����@�r��������
��dLeWp ���� 6���+�H.�Y7������M
�(׆�FDvfn�Y�����0��2�Xr�/�Wr����l�q���G��Y%}��������S��Ɓ��p��J-SM
l ��eYx���%(=�����b���c�"9�HlU/�8nxў"�-�igi�!��^��~��מ�%�eAhZ�e��omen��t�L��O�)��Ә0����ªO�ݞ��� �m�j1���-j���=���.Ҷ����$ѷI'��|z�UݤR!$L���ɤb�u�66S@�׹��3��ť)�8�xG�`N��(W�[dg*�WD�Rc��i9o����.�Ea��,��Cᙋ4��3���UOl����F�u��N�[|!I��I?���Bqۣҥa�B�a�Op�2\p31�o���n�����s1���^B�%g�"�������Nq}�KȔEճ�b\E�~����XA�!��e��P����8l�airٿ�~׭i3R���)�w�q���5�ê�3�('�G�d��o��Y z��e���
E�=J����',�߸�b� �t�'
��w�ɏ\�9����#�Ϳ;�W=ۑ��`���ށ�� e�ߕ���Q����jhE�!��w��T[H�D��Y��'9���a�D��>�Q��X�vv�������4b��v���In1XJ��Q�,HFlbR:%��:Qd��n��yNaѧ����p�<@�8Z��0���q��h7�:�'G/e�^��?F�	��.�V���>��yky.�M��+��a�-��W_Ñ����m��=�%Q�!�n��aqpB@�1����Wx.&O���l��R+���Nu�|uf%��|t��&$Q�_R+�P����3�99JL!ㆴ���/J�n�W��;�8'S�VB�]&�<,�j�S������D�m!U� \�'`)ޗ��C~�C�%HE��n�w�}h3C]����G"��8���VW�4���I)*���I���c�����7��75) i�u'{�i�be#�ɻ^�.|��[�Vʜ�?d�j\s �/�����I��>xW0e@Y��:�A�����cc��zQ��#�2l�̒n����t��6�$����Z�u��ݺ���w�Ɩ������N���](h:�m��2����,`'��p�����w�����V��k"i<��,I�����q�޶�~�����~v�ļ.do?��iz��g�F� h�t|P�L�cw�P�'�%���S�c�|W����e=����R�N�<V�U�����wDs$�������Qj�]�\�{!�	�E��h� �n9m��'����#6�] �zN7�4��̗
�Ow���-f&}�)��֗[�����{'��),�]��	�sh�NB�y����(��"}UP�v�~�s��5Z$Ѝ���9��j�.�U<�=�\���#��ӹ�/ �/ou�U�4���Ix:����{��j�(���`�~��T?5�U|��Y�o!JC�?/"�����`W�f%/:x[�`��~��c����~����!�g�J��p~�ͫIK�#��0�t�uP�C��07x�2�*'<�؀;.7��]|}B:���q?�!�_Vg��� ev,����2�V�a����u�b���6�ʏ����DDd"XQ���t���3k��"� C���O$dI��z��y�u��:�$)/$�6�A|
"T0�e`�[��je������u��'����K�q���ISDF��K1 }G��"�)��`�e9�:Dd��Eh���-���U����~�MJ!�)���ab\P�[H�"�D�u��%]�/O}� )�O�]�i#�E,�ciw�u"p%/�̰��}�;����c%�m�ч�{⪤�1���'������4\�̷˛{X��]�!D�RG��l1&�[U�`��f[)�3֢�x*7b�t�:Q�9��N[;0��N��/��QfP���u.QF^����5:��u�D�;���H\|��H����K�Y��<�X5�:������q&N�'���	��̗2Z׵z�,l�L�G[��_��ִ�jX����@e9�Cߞ�$`�d�^��.�K�$@W�RG\qѥ�n���Hp�(��e-�_���~�G�*��R�Fq	i��t&r�_��~�v�6����o/�Q�=Ҫ�y��)�km���v+{��R������=�����{���4��`���B�����>��
҈E�ܘ�
)h-0�����k#�Y��;[���*��m�ы�)F�V�4��)^�r��Z|;+��U���qn�Q��2BN�9�������{�-�!ҭ4�(�p�w9`��P�Y�֟�Y;�)<|]���T�E aN�hvaC?oMY�6R[��Rة�<��y�R���Ⱥ�n��Z������M�hs+p4j�
���Du��^E\�~���ŕM^S>��\����W���"�I���r<�ۨ�P�~H��*Q�C��ȭ5�A�����Q���~�N�;H����lor�h/�!��z���YW��- 利,���}*�)�f���h��P߾�
�bRpnU(�G��̣b!Qn��#F�"���r�-}�>#���fz��.�iΌ�ZP�2n�4�lQ����q�Y��5����L4�Nկ�\=u�yI�9�Q�g���������יʈ�Ygw��~�bh�TGm�j(��k')����=�y)�`�f&�퐆��x�ٯ� RH�$e_����l�����*Te��I4Rπs*�0T4G��\�>��91t��P�A��7a-y�Ʃ{����m�I$��x���� j�h����CJ*��ݦ�gT٨�"����/��SO)��'�+�\kr`u$�����9X�OM�y�龫�Ҕ�Kv���qφe+�n^1��߈���*���|)^�m��N�֓4�Ĭ�&�5ޭ��7=P�_�j}^����o��\Hy0���:������t!q�����0am�>���JAj`A�+A�����f�5����r,�̌U�G�\>(j��)�����6%����K-'����\0o��=�Cr����"��4���<I؊]`#�-O-�����RA�Z�Ɛ*t�!�u�?޺U�'j�a[t��B�kt�]�8�����>���\����"9n��34s����?�U�F9;�.�w����
=�e������Y��G�I������;�� �J���Wl�7�HL�s�G'�h�ȯ�,��O�A'Az�d^����L�ͨ#PK��07�75b An��H�Y������<�yO��s�vC�O��G7r�d_ᢟ�f�ZQ�ɽ$����� ��D;-����� �1��o m�9�xͬ+�
���+����(��:�b0�w9���aoy�"��Y�qdh�1'mz�f3�Sey��?���y�יT���W(��f����a��X��,L;��o	
�����*Rκ�˻vLڍi)&W�:-H�(��i��:1�j����&��"��Q��n��0������M����})�y(�t���bx��7O��'�{�Oܛ�PءY�%����8����XcK��!V&]�5rk���@.EYΑ�v��YY��f+E�>V��~ �U17uu�n���Or[�y�X��R��3�-�P�Υ2�Ǔ^�%*3�>�>Q�Z �]@%M�҇P������}�xK�A�T����%N>4��y�C7c5�S^6*�r�`�(vU�QQ�m����_�6�\'ͥI98w�T�e~���Z$^��ep���`��
�R��v�7�D�s�x�$`o�,��zb�RYX߃��P&RG� oN����n�^��V��~�Z�����}a�yEy�)��y�N�3�|��0�ڊR����x���1.E;�$�EV1��H�fV�|�a`g��m8]%�3Y�֗p5��4W?71��W�yE���� f���(��	B��,���f��ҹȒ���3��a�$�/�Ѩ���a��X)��I��L�T�`&{Fi�v��:v���p���4��R����8�Y�����:Iмy��X|�wP�A(6aQ�T�q����x��&3XT��u�'�q�|�}ݡ�}Uk��#Y��dF�l%�Q ���$�5�*!�����KT��#��D=0���N���(fw~�����]�G��7�I~歐����N�eb�gQ�10�01m� ��-��G�*��RČ&O��+��4|���1w~g~�ț�2Z��͍rt����/���.o̸kh�o�K�cz^GC�o4�D�T�>z��N��G���	�����14����KK��bz�G�bL%��3�|g���-�b�r���*��h������L�'�S	�� ��g�P+����ٰ}Y����cD(��Oٟ��)�-���ࣤF�z C ��m��Q���&k�&T�Ԁ�sC�"�*��R.		���O�Z�˻iݝ�-C�p��9"QqvŜ��9������� ��5S/�������rof�+Z�P�4oK|��K1 )����li>}�l'��q�+z���y�3�������ߺ P\ �-	T�@�N|�ە�௱3����B���6�C�9Ѹ��l�LT#+K���H�ØuI�rfW�zA�}2������}i@޺�܌o�����)hX��u�(\Ř�4�;�� �	cg����Ŗ�����u��14)e.l�Gk�2lY��d����IqO�z$��C�	�S���A�MqgWN��Y����0�:���7�m!��S�"z˘�S���Yŭ�u��]�I�<�kz���~�"�CK���2���_��bvE�6>�bJ��#k����7
_P耋�{�[j���S��8"ҨH����Q����rms���h��u[�Z�t5��R���.�F���2U �O�,P���5�2�ƯX����0L�E*��������˫��k<P��}�����|Z�z����ړ^������B����x��]�%ꌪ���o�FJ�sp>5o�Kn�]�ǳc�4Ԭ��R�Y\6{�0��")�X�%��g?�u��(��3_�pKຌS��t��f��@�=����M3:�]�hQ��oߴ���ԁ���%�+�	����_�%���}B���KU�=��}�w�Z3�=�����hU*,�>}~	cU#H�cn��ۉUԳ�;��\lv&� ���`3MԂyUvڦiaa��� ���21v�_A5VI���*��M�x��F�_..�Ecl����i�3;��H]R.��ho�\?�
^*����1���up��rcH�sZQR"5j��8��H-�H���Yv9��ylR.[q�<5i��$e9���H�_�2 �sJ�ß`�k����>|��W&(؋��/�[3}���@��;�}��M�+�����B���!��2���Q�JU ����i�b�@v�'��4$͡��Yi�L_^0s�ug�?����\Xz�4!���)�*'uGY�ΪYAH�$ݓ��<-C�jCVE���9#αE�53�R7[�J�r��\Rb=O\�����Z��z���r����F/�،g Lx�D��(�eB&	��T��	#6�O:����:�YT�o�W�hB'����$�2V¼&�b����N���v_�򚍻��i�� ZY�������:�表3nw��3\f°>�4� i�<A��1v3Aa�Z�=A��n��i��e�|�Zcvx�·T���
��r�{c[Ϫ̱�L4��gQ�+Y�����v�Ҡ	ݏ�G�8fR��NZk��%�����2�Q��`v��m���H�b���E��[.�[!�څ�L�lu ��רK�C!%�z)��"v�_L���/��/oδE�!�[�L���_�!���(�� �V��-����G��ͬ�� �TԢ���k��n�4MX�N`�ߞ^���;"|-\A�W���vɒ+���WX�^��;�x�~�e9M"�@.�������Q���Rh=�WH���'4옡k��4���=�x�8�`){�����fl��7K$0��Q���~<���Xn�A���(���'W��r�'��V�[3��dQ'�)�TnU��ƅ���l�?��
��I���S;/�\/+ʴF��3X��E�9Xuqw����g�|?��٧��Z��J���lJ�u�5�@4�Յ��>�	��zs������JZbP��*_�˰��Y�}?
,��������k�o�0l��ȍ�S�'��?y=D� s�mӍ��S�����O��d�@��{����������B�h�`��}�����#�G�cx���`'0����g�#�J�	)D��yA:����)/��_�n�O)��q3=���	�
9��έ�e�;Q��V`���:?l�q�G�s�İa�yJr���5�:&<w��9:�&�g�6��b}Y�@��O׿f�%���=�9���z�{�nشHZ���#[��B���7�)i�t77��s��닕UaB��+�P����G��gD�%�ҭ�F��e*Gn��������$���ψ�+�����^��e"I���ל��>E6Hù�:�t�����L���|��M���|o���y����A���pE1{�Ըِ���	;�����.��g���G�P�K@U�+	�k�K����TK ��]sC�ً+�SE�Y�75�a��Pk��$���c�5�R<	?��c+�7�#2��XFV�����bc����ws=V��BoS�zQ��3=�sn�.l�,bTV�4>�A��i��\���Qg��9�c��h_��v�a�mX�-�� ���e�̞T�C�하*A"�X}!�3�����Q�{����'�;�f+'
��%I�"��15��߱��!����;����Aʨ�j�*���^kT�jĠ�+��%V�w��$��-QA�3���Q��m|��ng��ĸ��BM���E���b�"c�X,�����6��>�=_�h�R�܄.���=9;����=؄�1���0���b���Mv�n)b�����+�I���v�g�Uu�!ge6�BTT��PI�5��5�ASB�?d9��C��S�%F�`�#�A壇ZK@�f�`�����G����Fz�|�v�%x��p(a��&4F$f�پ��bM����`u�z���&����T=t�����6��_	��&�2A�	�Y�.ټ儰F/9;G�r�C'��"��PAcw�����xr�0��2�����B&���`��A�]`�a��0�++Kwо��o�d��e�6��~�L�n��Դ� �x��W�·l��E�E�57u[B���q[�V&�Mì��f��ݻ��]��$���?���A���|�I�煻`�"�}���p��T�p9,����8�,o"5rxZ��4L�)͡�W���\^-˅=�J':��$!SQ��O�0���P=�\�n�q)���:�Np�����j�x�7!�D[�I�趃�f5il���qi?�1s�;��	W��H����tU$&�����=�RTP���O�zxto�� ��7���w�(�vȝ4�#���q���Zot^����Ź2�0�[��ަR�|*U=ߡ��~��H���\�����j�0c�d�D��j�HTDP}����5$��,�g����#�.���0\��:����(9'�F�ٲ)�0�Bb�n\YU�E�M��v��Q�%����`�������1֕�L@�&I8��AfǀJ�g�1��܇�:�K*���XuRY�Î�qt6�U����x|��?��� IFWN���
(���DU�.b�+�p�O�a�+v۷\l�Mo�����I!� �|�p~e�3�#@Ԉ��x;�� U*r�m8��p����N�!d���¨q�EP�����F������8�d���o�H�30:L��:�Vr��&)�],t�7�\aV�U #:������m&1�N�=v"j_�M��2+D�F0Fޘ����	�T�Ug���T�/��X�t�]�PR�n�ELB8c�*q�m~{;,��O�MI�5b����%��p��q{�+8`$f��'�O��1`��� ��{ָ1l�{t�/����r�3�$���Y�c�x�[��^LC���*?MX;A��O����;�R�cVݒ�� ���Cu��n��R�;Ew��'�u�<�%:%�����Eʹ'�t-� [��dļ��i���]*��z;#�h�I�Au���Xj���L����d�0���)X��Fr<&,��;��rq�x$�2�k'���G%��BiT��	,z=� �.�	mf�;=��)��y�0���Pg&����,�H?	��������ugB4�ˏ.u��Do���|�zD}��$�7��)�̄y΋�"��.*�w��9R~+��Ub9>����xb����b�ͽ���G���ĻR=�h�l\�l_�EX���y���|3�Yi,��٩�+����<�0�B��]l��: ����y���w�y�rj낂��63����-̔�dk�EᶠZ�R�D��t �����a�N�Y��$1�f2��s)���Q�(�o9�N�N�d"�<�:�����'�P�i�
��W�z{�HO-�}���3�K�p�|�1����nU��+��~�*5^�5~��QAҌ=��h��JGX����\y��Z'��);�"p�ƒ�,�� {UP��)V�q�U��y�Ft�[�uy͎rUm���PV	dl�ӕq�<�{� HH';!Z�}$��_��"Hvy?@K�WY�h��|Ơ��,a��?8���NX��ڹ�	:��]���.RXZ��T��df31����%[>�V0��i�$zyM{�o���yت�Ž	���e���1`}Paluϲ4<~A�\�Mj���O����h�����	o�o�z����=�+y�	���`"����sش��p_ȦD��E�Z��BA�"B�#����L�He����t��C��չ�=P�Um��a[��f�ì�ySS9�M{1s�j���+wt������ۘ�A����f�,2"Z��vO�v��5���3i݉Lм:k�ڳ�ȭ��ؒ7~�GC��n#��Z6���Bt���%�	ЏY��Ǟj����^2\���?G��Sx�G��5E��6C7~7� 0N�~����;Rg���E���+nj��׋FkX����Dmq��&,�t[g�0��=��WoEsVP���gV&\h*҃q��!0�|xn�iO�N&�;��� ��S��g0 �6��L��SB2��&޵�y0�/�p��lNrL��0A��Ҩ�je��	���]�L�-e���E�[�,ہ�2�8�K%J8����S��@��t�3d�f,�=�FPym��R�x�p��h(���Ou�`��Wm|�O�wz0Yd��?��M�o_�k�$�Y�+呆i�d�ء�x҅��q�M�N�_
]�D} �Nf���3W�Se�4��D�.wLAd���h('Kf��_���sxߡ�嬺�6�����X�B�ur�c�n�l�C��������%ϿӨ�Pv_.UTm��ۂ#��ϔJ!"�/����//�6�ߘ�g0�ߋ��XmR�։u:t�|x����UF����Q'��a�'���tC�b�@�~2H�4���(��ۢ��w�Ϥ�7���pA���p�k8��M�
bA����T�ؓ�'��l��eZv��:��>�R�����V�;�R� ����E!�ۿe��S���]��v���Y 5�d��7w�#S,k���n�Y;@��/�#�9��f(Ge�F�h��T���}��|F�T]0�j�U��0��z��(	���ن��[2�%	��7�ⱨmXvwVs^�U�0�\��ـ�V�	��u���+�Oiw���|W�V��v^P��בb�)YqX�JW'�qB�q����P j"WO�����_��$L�%��n�f�������'2�w��|�1T�M�B�������-B��K�0g���ā���8�1[��m�T���fV���~KR7:�;�E;�Ds��9���������U<�Sj�}��A�AGM�s�D�r7!#X���m�f`���$M��7�:�E��A�)�!�R��8Q�V�A���f\�1n2Z������4�%��|_}��D�(#kH^���e���cH��.>&T�z[;b"r��6���C�)��ݜ3��@s�dZ�G�eѡ侤�JH�L�`&J�կˇ1��S?�r1n��O��GU+z���<�АPTE
�g�~FF9^ c��{��f�i�[A����H��ooIVFE�Z�0�瘛z����yg�����>� 9�{"H=� L��Y�Tv����ix׶'�<���	t�Н��-~�/N�_�cł�w��C�l@\��k^2�k83�����Gm4����uk-�����ֿ�g�b���.�%"-��Rl4��pO���F:���ԩ`�iS�/m���Q�V��NĒ��!&S���y�j���o�D�;9%��	�~�KOB&��j�Ͽ�
�N�����Yr~֊�e�m�K%�w������GC�L;�-�'G�6�8t���Gl-��4�2E.���U0� u/y��"=%�S�mfh%�Vq�?�(����C��G�ϭ�jy���0���p�?����&�.�55���U<�[=H�c�X���bs����w0D�I��I/F�p�7/|�}�#�&���mĘEfE�8���ۢE�n����Q���i_���Z�c����M��fV���u�EP�]�U�\��,d�Q������_�\�Xn���gcsk�'zRw�.�A���#�%��Z�2.��,�i'.�����ړ2�%�E��lIc��;���\6�1�������M]��ইP]{����}�f�i�Xt~�#�m�*o�X�<�I�	��\�y�B�,���z��<�(�h!�u��Ј�����3yi?bx~\R.�[�7���l1gp�ڄ k�P�J���Dt�ex��śe^��6�fn��H9W���ք��bXLc���Rx�]|��,�a^��¾K9(��p�'�0����%<b�;�2Is49�P#l�We/���3י����֧pƎg*]ϭ8��^���#���O��h����^m�q���d�:V겱�K�Z>P����'
F�}W]�}Ҧ�7"�帳@��	�ı�)�;�Z?G>n ���N�e���u�c�̻H2�V�w$r�j�]־�۽C�G�_ql3F)��}q����(���:�p�m8�Ű弑���ȃn��t��&��	w~�#=��m�at�SYV���,p�����������:uڼ�8aw#H�[��pNh@p�S�Pz��ڼ#�j�u�~s�@�e�~�c�	 �4�X�����ㄏ�ک��k{z� ���\�f�G�+;K�Y�'���W�%��ՙ�mc�ٟ�^�)�����)����XJW�J�2�ذ�kjJRy�v��t�UiԖj}��ּ�����j��!�`N���0�y�P�`pc�s�C6���`�B`Dp��R޼nW�����7����QÉ��W���1�
�f�?�ҌR�6�4M��4!����cXދ�"c�y�T�_^%�yۈVE	8�N���x�q�q�N�+�f qL.<�ħ�ԃ=ב�r��8|�7�]羃�Y�=w���mi�j�/�ԳD�:�/��M�˯����s�����s��Ӂt�(V�M;~���1鶼�,�%��f��3�kB�<��sS9YS��K��i�W�ѥ�q�H��F�UѶ�T.�=�X��D��]$�e���e���;+�6y����s͒>�y$�%�]���^���1Q)� 
�v�����E����i�;p�xH|��U��~�f,����&�a���.��]̦��6�QU�;Ll%N,[{�u�\��j	�D��9�R��NMY{<Ҽ/�U�� 8��F�
����W�x<���Q�i�}�˩������뿣%���T�օj,?4���n!��{|�ȱ�Vu�b�����������oP�OH��wg���ž���h�>�l'�8O~����!��?l&����ң|�Q�J%V�H�Kα&���B��������yG������6��uI��.��T�W�U�y���U�;��0{��c��%��W#�%K+���!���OR�S�����6��<tj��S&���:��[��L�1�������/�%����I�:v�X�%k��9�5�5��1�O����!�>3F��X�<�L��n}+Z�:���z"����2e�n��O���i�#>�0�X��f�K��vg�Kif�3.V����_�&�\S��ԛ�)T��#��3��Ć�iɊ(�B��@����U��o~�aiL򟯳�$u��HRx�r�hK����~WMnZ�R(p Mۋ��t @�gL�}G6����X�;����`��p�������.$���+��U���0s�9RL�e�&-w�G")�VU7`Ӄ��G;q��B�3�����G���uXG�FU!MJ�2r��|v�	�XK2d��(&�s�F'�3�[�L��<��╱בF"T���W�1Ad��W^�	;Y��i�!����P�i?���t�M)�֨ǥi��j��M���췞7��ss�	������͸�a���<�/�K9����R	/@�iJ�;��c�!Ӌ�.��$Xo� �z'-A�4�7�&	y�<$�L�4�er��q�9��i]��E�:N
�h�\%~�ݴh J�py��L!N��@q�yT���=�C�:�z�k�D�8L�vJ)�ܹ�BӺx�~�z?�Rn�tr
X��F1��D����(
��-�1W-��˽}�D嶵~|�ғ�5Q�����4Hɫ���R@��=�T.�O���
�c�(�7sDa��[�#9��9p��g�Vm��ZmF��W�����k7.�P���G�ܩ B�[h��ןTX��]|�g���5����ga��P�u�O&C��G��NF���K�����z?�S��Ռ�5�T��4.|t�Ԍ�G���hl�&xd��ɍ?p`�m���������ʛ�my0�펷m��8��6ֽ99�P���_IER��E��kߞ�v��5"$u��ͮ95e(�u���|9ܝ�BZg��?�I�E`b/�1�c?y�d�N���j�����TE��c���ϱk���.�P ���S�6�U33���@�)@��M��miB,
s�Y�~�
@)��UJ`iq�_y� G��
�ʽ��MO���\f�OM�]�����A������5�;���Z7½�7�B4G����)�
r���CM�vH�I�zJu�LQ(��u�Esc}d��^XE}�h����y�f���'�mK]�Ho�W��.=�_D���X�z���T���_t���1�7�G�+�eg��=6��^�� L���m��>|Y���u��>�p�,�B�%[u��[&H���kO!��k���$����]��!ɖPr!N�䒫����u��C�j�.R�M���1�L��Ԯ)�='?ʦ�>9,��� �/�4�"�+HQ&#@hؼ��Z��բTɈm�;
��AV-�̦E!�Ci����L����
z��:�E,Ћ%����!�ɞ�1��'� ˅��\��7�W�S�˂[T��S!N�ώ�U��cj%%6�S�
�@(�h�o]����<�[��i��xҢ|���_��ņ��YE��۞�ϯ�uYnao	��3�7�/�:��y;HW�_�4pL�^�n�!ԩZ�p5�Q��J�V�J�Q��~�5 �,%�}�QZ��2�R<Y{s���1�j�J��ε��%v�R�7�)Q'�ek5�nNJ0�w/����MnR����E�Gv���^��I�4*3�Xq;0{��8��׏6�4R6ͧO�Z(m�_)Q����jZ��\i�]�F���J�a|i��)u6�]���J��/�{f�;=�6AЄǬ�Z'�Lhv�:� $�/v�%�r�'.�Ӏ��Eu������W���V�%����#-�������ǕY����*�ɠ�0d@	ޟ��snc%d�W.tۛ�h,��������$��;r����D���u��)���h��9����=��א�h������C!��%=g\��Y�����4nؠnǃ��
�ϳK��Y��j[*SR�7G3(M�����T}��2��4&Xz�-)��NO�b��୛����� P�u����>�ayf�I��1@�T�C�Ɛٝ�����y������xʭ ڿ�	�RU>ыDfH��SQ�x)�g`ḓ��9�E�p�e{���C�3
a^WͽQ:���c.s�=�S��(r찤mO˩j|��n2���9����Y�r��}�q˔�Υ*���!�E�S��֡[�w)~��S�K�'ms�7]
La���:�G�ɫ5��zH�n#�<}�W�]'.����s��H�}�=�VI��EN~�N��{��ʦm��Ɨ1�V�!&:����n�O~*ی��u[SubX1�\2����{��
�.`$l���2�w��T�GBgs2��Y�'ATi�S��A�㱝1�;�u��9�c���Sᩲ|h��|��A�=��=@Nσ���`Aw�^zG��Ζ�}:[ ���p먞��
(1Q��a!��\c�^��9@SZ�Ĝ���7�Y>��x岟���I0$��p��Y�k:>i��[G.�+@_�uV�^k"A]�Ρ�����_��S<��!!F�+g���M+�3��POP援[��O8����33��A)�9Sk<\֯��>��'�XI8�%"żfn/2�ϰkJ|~�����s��2����Ҝ٬l��e��I�f��@��ڵ�l%��$eװh�,h�8�R�[˚�H)�aҝ�e+�]��ˮf�s�X���K(ֽP�4�&x�|������*8���Q��ʰ:�H
N�i���0 �,K�F7<�Q5�$dT�x5C;��äb�(s�Ec�w��M�e��[����(��E��q7�pG�xN�L����My�hQ�:�(�WKiJ|d�	�\b@�dvFX��yF�C!�c��%~���O�ϑNtu��Z�]��4���Qg�g�g�����gS����^�̱Ʃc!�$|N�Vk3����s�l^�+p%�{�R�1��L?��� ��6e�2��P&Y>z����IC.B
e��σ	1W�}�7��k���[;��;�f�N������SW�ʼ�xo,P{!N[�u���N��Ra�l;]���"�ć�u��`��<���Un 1��te���M���)�$�٧����@���������p�5R²y	*���U#.{ ���r�;*�[D��h;IDb9�F�����i��t c�K�����{?����ѯX�b��I4"3�;��A�SJ��@������}�Ʈ�H�3i���h5��>j�w�mJ1�����c�*��G#|@�%Pba�2� �]oN'��0�t�m����s���q�X@ҋ��ӟ�����cT�>��\4�cD���׮�0tHmW6'q�\�@��ՄKήR����c���x�)N��m�������5１�d�O9���{�}�J��Ұ���b�4ׂ�L3.��<���.5����!\�Љ��A/H�#�jMu�f}����N�\f@/��pY
�7FY�.>�k�{Q#%�b�����xI�.k "�����L|G�	��Ӌ0�}N�r ���8J�N߯����uA^5�^9R?�-D�i-t��m�|������[�B_٘�����U����[�Bt2���C/��	�L�|�#x[��Ju��V��GE�8ky0�R��-
��{m�|��/�>������)Wj4�^7���[r�Io�cK�q1<f{��;P��^
nN��1�_15�3�%��E״%W)�@�pNo-�d*tV�`qU��q=��		�ՙjΈL"�Ћ1^0����	~���v%:��ra�}Ss�l�f�ܙDA� a�9��梥&^����+Q�7�����:x�2�kK��;>֯%����jZ�TY�6�1	�cᝊ-C�j�	n�e����x���G4kT�@@yT���G�v-�E�^$[��r���q;	��Q���=�I�CY���V��D��_��읻�j��?1X����|��b��t��d�l�t��&-'�-�5;TB�p,JGOw yx�w�L9v��'�@0ى(yY�hb4+�7�%w�|��ɂS4j�C< ��F#2ǵ=yy"��w,����;S��Fњ+Jo-=����Ҽ��EluHUZcE�b ��z����h�w�ݭD. �ީYz pE H5k��"n�l��@vA��{+�q��Ȣ��x�{Z�k���r��/"��5h**��>D���7��g��}�,�Q�����^�
�+0]�N��w������:*�R�A��9&8��k�+�vک�I�h_㰭k(��)���%��/.�x��8?״�_�I&+և3I�v��v=C�VU�s����S�21�����%$��,7V"q$iΝힶ�/��~&0}��P֍_<��<�xB��o�����=�u������c������

he/*w������k�S���MNO����P.���_��u��Eձ�NV��y�'q�>w�+������=T� 1����n}���z�5h-ޝNܰNy�@}�i��D���B�u����d4�]�š�),�Ͳ��Ĺ�c���y�Br�GՎBگ�Ŭ}�Hl�$΃1.��ڌ!�8���FVƙq�k�?w���3KdZV�r�\�&���X����� �Ur�x]3�)<n�ܬG�e�:F��#4�M��3s;��\��YxhR�?j�U!KJ�q�|
�
+ ���P�zT@*��
$���66����K�J�9(���Ȧ\�	�a0�Sg�>,�J,@q�{p�=��&��L_�{N�\�� R�����(
*l�v����4(�B6=漢aвW53'=D�@�.]�E&0������U��X8�6W�w��{��� ���(��A���΢X/LƩZn�N)���pf�P����!/�+D+��E��Z��!3�
0 �~F׼������O���E}�׊f�]ڹ^F5|���w_]��l��4 �e[�e6|��#������s:4z�o}�Qn�3�i�+�hn�l�o���tW�� fF�$�_Fʲ���KsX�9�^�L F[OS^�2j�N�r��QJ7\Ϯ�ྙ?z�R�9�U��Sp���o��eQ}LE4~9u�|]nP#q�$�j����B�SY�pUO�Pr��r�.�}P���Jɰ�ҩ\�l�enZ�¦�T�~?��+�V�&JtpwdI�DE� o��0e��"aѐ���`�e��@I��c���ĩ�Ig����dQ`�C�^Gc���o���aDo](�^�F`L�w���L%��i�6=1!yU@7K���s���	r���%�PG��]6i�����ꎃ1B�� ��������M�ˣ�,��Ҥ6ˎ1R�٬T�vT�-�$u�'�u.�� @�[2���G�o�݆�fOƳ�������8��s��7f6��+ҫ������V7,�WA��,h����y��4�����nl�A`��'*ϑC��s���[�3}-��3�w��3;�����2�X�%}�wXGNXp��q�E>� ��]ʌ*Fu�,�Z��l4�Hb���{�|�S��dT7�[����K�����B�mh8Y�pl�63)H:t���� {�y�C̑Ȝ!w�~T���S)R���/����(@�'/̖��,
Ic�,�fJ���S�dDPy(�3�y�c�JC��lZ� E��#����"4��!9�)��Ǔ�>��q-D�ps�:[����F�����'��B��.x�nvaߚ'�	�Aq���[�K�;۠��}PI�r�b����o��m�膆3H0El��x�"�K�����*�Ĥ1P�H�:_�[�-niE����m�o��SNf�K�&l4���|^�D�{�f�~�7�"�L>�
x�%���dTSƟ��yۉ��hu8�-�-�������NA٥�6��V�?V�S��1VX��f��S4?�7��Y��uLg7�m�ϖe˘c��[&�� De�0%�ooI���o�%�Q��:�j�m����+CV�/���)������"C�;�p�zEP}}j�)�����B?n�1���Y��M�����C��*���Ba����2��@���0�ă�cw�xW��Z �_"�Z��=��Zn��̖�� �ʩ�`�S��s,�v	%��D��y5��L7STk[ծ>B׹�R���"��KF���n�I�p	��͘`9ro��!�W����� 1�?����E4��?��1�JKRI�?��	�bd�7�6�V=)�ԋ�(���f��P�sѽ���x|Dr�[��V�1�^��jU2�\��A�4�[��H�G�5����R-ۯ�给�u���D��p݈\�0���:�˕L;��BD�I룧i�eӓz�$m���������R������R�ڌ����#��V�7�W�d��[�� �e6�S�S�{� p��s��d�I��i�$4���؜)�[Fd��9ZP`�\��ᆴ��*�P�%3�C�a��%�q��H!%]{�������2���X���,%K&ߍ�X}W��B�g��L_�O!bF{9���h�^�4��0��%��Ŗ�a�?c���F�d<�����tR~�nA��t�:��p��1�XlB~�Bn�R�Հ���N�Ys7&,����Q���NE合�YK�%p�L=��x������ /������sO�Fz�Cf�,p���Y�7���kߵ��6�����?�aZ΋_�rG���H�DT����a�vz�Z�	�����g��7�b�E��.m���q4uyHTJG{˝���c�"���M����W
�xh�g�d�(qD��z��N�I�c��'��H�t�N�����UT#���LﳷNi�6]�%�tёƶpGɊ������iyw��U���=Ie*�+��S�$�ڧK_����)�>�ə3��$L��@�- f������g�ꗖ�/u(���~y�~=����ܓ��PUy?�� L0�/�t	`R�U��+�5?c0�.i6tv���O��{�;��,�K9�7��JIhI��Q�Ygp^��ء�B�>�[`ri�9�����s�X�p��cX�ϓH(�r�T��ua`�"�f�251뢒<2K��~���:��!�q��ǲ��bt���1������y\��s��n���io8�$+.�h�l`XH��?�"�����[\��@��ǈ��/gɹ��`���S �����1�{��sX���‷�ܸ�\;��W M�l�o+!��b��/�Mv��l���v�N�jo�%�d)�Sڑ]*���?���G��D��S���e7-)F|��Ѿ�,9�Zt��x$k�A��ٷ׊{�������c�Yjb��۰%�%³�܌}�"��q7z�Ê��<ڪǡ-t��/6U���Ӗ��sn��[��c+��o���6�Jx��K����i���V�f��$9%�1�zID�C O d��su�Sc"����B�ə��ہ�r�x(�L��\Ȗ�¯e�լЕ�,��&u�o@�!�'?ﮈ�<J��_�x�ڳ|1��݈�� b�2b�e�hg?�t���g����ޮ��ճh홭C�*�#��ڢ����N��8����,S^�4��w7�7ђ�=f���C�g�|7r��ؖ���LD���U_Er�6-׸Ы��S2��ӆ�[�S<&Z���	���B|�!-w@����7�f���mM#�(��">kR�+�c�hgv�(-�Nӣ=�+����н�eeAM��,.� �ص;H ��K��@Ja��v�
�����u&+�S��r
9�; H���ֻy%Xx?��	S�a�P<�x"�P�	�8��ڴw���h�oSN�z�tyg^�����!���'��L�_�/)?�ؓ����n���O�>Y����_�]�������Z��e��p������d��]tfFAN��n\��Z6�#]*E��������^@"�A%UM��{B��L��b ���l�%y"n;����`��*5�7�,�a�۾���GPl_p~_U���g��(/����;�*�>����Ut�7�^�HN^��7�2�ً��~!f9ë́H��H��:T�i�Z�˃ �����5�,�{c�*�\�PWH���O2%�B���^�>=KH�==��M�|{wN��Z��D��r�����H0���+�&��mАߙ�p�~b��D�O��t��t9[�6���#߇b06�w���0���n-Y>k<mx��Z���Q�-���k��Q����Y� ���*����㊥��X]0���h�=��Р�t5�H�u�C�r�_����;��u�y�qlBa(���T9g��87����S	�-�����w$��r�<��S[;�eG$�*K�r;^�q0\�4�h���Mz�����ޢ��64���d�"c�-X]R��5}��D����ޅ
������~hWH/oͨ<\��R�'���Yv*@EG�b:A��}��*i,�������ϵ���"ܻ�.����F����Ah/��Y?\e�Ѫ^��Ԣ�C�� &�AΎR��h^ee�JXA��
lw�a��!X�z�NKZQ�R�Y�TDH���3U�U�KK�Ʈ#�nՒb�� ��G|�<�yc^���4���I�p�T.�1[\ր���^-��A���!鐒���x͚bZv٨�[��H={.�RM�U'�������H�s�9h��`ϩ���Czv#�Gf�:�ٯ8�s�,�3��	|/���d\�0�=���� ����g���]������O��R��F��N���vo-�b��=�8*oW�(�Ϯb��g�TXr3���l ߪ�	�٪"����Cݍ�*������C�� ]���T.dx}:E#��'r���`����Z��p{Y)�|en��T��J|�-�e�G�`�l����DN�򊟳A,��]?��}&�2��hQ���%ҝ���wd�'2��[�xEoo��F� [���%�� �`X��Ƅ�[��D���/��PyrW�v���:������iT_���Q�'%�b9��],�1`��ǫ���cjdlw���D��~F ��J�zPq0/��~��t����e��3	�U��lv*�*��v�A"��r%{+�l|bu���, �_�5[�93l��0��å5R��	Љ�0���S�]���ښ[�4�D����(O�� Khfs��HuH�E'΁>�L�k��/���Z%���ؼ�
���7��Ie�ja���"RM��<M2�sՕHP����X� ��U���;��k�)}�l��B����l��s �oǜ��:�J.X؀P��L�G1�:T�(L9>�3����?�ͻ58SW=�A
��ƺG�*�AT���"��3�O��҂L�Nj%��t�a��IAc3�&kюP��p��{�Vt�ץ �+���/^q����./��&�>���Lr�����[��A�x��Ρ*޶>�n0������a�5��/�
p�y%� :|{T����b2�SD�UrF��چ�g�٫L�|�߆�$J��w\ҧ�b����_l�pק]g��'�n{����ؐ�K��\(��<�apz����S��_�RD��~(�C�k�4<ƮHk���m6��.��E]��45H�+��p�^��������?62�|�A0,�}�K*qL);�E�(�f��(�`��Ӝ.-�z)��N���&4�]�@�|3j��Kqk��?�0��p�5��x�P'!��v�����ݦ��2��N�6#v�G��V�c�֘"�c\5q枮(�/;yw�Ը�(
��C���T�Tnl���!M�iCG1I?�6�+e5���$�ìJ�_�Y�!������E�)%�	�@WT�������Y_��
���dtH���.ȱ��գ��ߣ~���� �R} �t�����%�/�T��unSI'�W���)��1�Xr��%�2������hQ?�!����W �?b��
�$F-��C����j���M�\�� ����'w��R�өHFrc�O�W��s\I�;ߧ���aO��B]1�(�i+��!-�	~�` )E ���|�|�SE��k�8im��~�h7��k��w]�;�޻��9空��X�/)ڡ�g�I5�Wh0�8�FҚ���H�ol|}��/��)'�l�&�Y%�u��
nh�s&_�8\#����h��O�X�Z�������s��I'�C*&���}��>ʶ��tS�T��ɰ�g�A`�\X�-B��)�� ��so�'rLD9̖l�-ǤoZ ��j�����af^�[�3�9��Ms�ȇC�J��5V|��@�:IL��	�L�%�u*+8��G�;"����A�ؚ�B�9d����hM��Sq�}��?�ޚ���ױ�CxH�>����i��L1T���I�&+x^-�D��`��*4��^'�q@*j�Z�"-	���͜�6�����i�P���+�����6a��y���L�eD�7xm%�e��D���eFB�>��:kJRҜ�`�ڌ)S��x�Dm�>�z:�v7_�2�]����MH]`
����A�J��+s[T�F��c��JH"�Z�9i&�j�$��s�������s5Ǩ|��pȜ5��G�ۼ�sW�6!�S�	���x���:G�n���zQ|y�>�s�):��_�Lַ��3�i�!�0���T����(���'v�KYPC����b���y7�M�4ԥ" �Q|>�'�<��F����9��߽�[�`y�bƈ��}�=~𬙻�Oi�π����Oвj����r���9�u�x���͌��0��M*V>M�(>\t$�D����Y�B���+�7�����E:�1�n�������
����{;(N��sJ�Ms>e�B_��"��2@����HQ������]R��-��?�:2�0���wk=�z�8��PXZ�2���.�Ð8�uu6���~�dJBػ�+|����^c�i�0u�G�ɏ�ʅd���^���Xj�2�,��ŵ�k��Ppѥ��g�t���	 �T�P��3V�%�h�;����E��kj� ��P�hT�����uŐW�ԝ����'�����;hb�2m�6"��q���|$�d
��xs�Hm�뺾rA,7�`T������C����⼗��7@C�ׇd�GJ2��P��/Bt��x:�0l~�|��z�-a�A.���Ի�h<8�;���tR<&�բ>㘝��F�O���u��%�\+���V[EaA�NET�.��=,XNi��,E^�����陈��JEJ癫@��%�K	�j�T�ҶW�^T�ʲ7�͜�����~��N�Q�B��T.���ǆ-i��6Œ�`t4���|�Qm�������X}��y@�=�6\�-&wq3#��Ӹ���ǯ�AI���gok��e+���1�;[���>�1|N�>��`�]6�!d�Kyp���\KpϣUo�])������UV����ꕞQ*�%��\CF���F��L���C�V{R�xv��ai�G9��_Yº�J��.�:�H�\�SF�I���H�e���U�
�iI�t��F�E�G�^Z
_���Wv����l�������{k����{�vg�����E���#�E(��oi��B���L�㺇J-H�X�KD�
�P�����%҈��\tbR���K>��=���Ee�d	�lĒp)b����/����K���W7�6��$}	�:
��N�S�*��e��2iI��*�wFtM+o���w0��k(	���M��g�٘� ���[x2�Ǟ2[��H'%y�c]�>�l��C���]>��Q^�=$6�/��s�C:�p�,ma��GG&D���m�S@�Hڻ�n��8�&��f���X�~��C_�l6\�G*���}�`&�vÂFtu֬�6^���]����&ߍ&�;>U��Z�,��!���pR�&��VM���� �e�������Ǳ<���[']��w:|G�c��{:����^�P79��ꄀƇ��Aj�zj��S��V�ET�Z_0��Eqnq`��r��)���	2�[�;��j�G�����6|���ll�ش|7�9p;ae`�#�&�kY����0X����h-Pq�,� �'�`���n�W��J��)zȅ�/Wb����γ���>�$���c����Wb��9׉<�R���B��2ڈ�:�o�I�4K,��[Mgf� {'$��.	g[�J>�	��sG��+�����(`��W�/"Tj$�"6�T| �E8-J7��%3Dc��7g9�2y'B̈�L�X���K^��D�,Q�eCk���ȝqK�u�=݇�2�dZ�r\A�P5b&I ����NC�	�f�/WD�6�*o�o8�gXb�xylW��%Aή�z����T�`#?��=0�~��f~��Hjw����e�XC!��/�6�n���Ȉ�t�������|z�b�D�To��f�����賾�rAΎ��n���2{4�)��FE��їmi���G�*�%	��� vQ��
�~A֑��f2	&A�3�3�JOI��ۏ1��I��UҽB��u�2�^S���_7B�x�����k*��>J�6�5�헻Ե��ݶ�~�.5r!����n�`�M���ӓNy�� �5�'��l���؈�o�ӣ�`f~��m3�;��p��O�G�7��k,�x�i����ř�(�9��XfZ/m ��G*v7ɽ�����\h�wh(|'?/� /qt��lz|��ֽ�L�B Xg
x" �����'�7�8�PCK��/k��A��M�ƨ%���#��R�#ƞ�C	L��=&B"�,!�-.�e�g�]!;��a�^�)����͆<�0����ϙ�A�����<�5�#((w�Qv5_�cQ�k7����͘*��'�Q���bcL3h��etݝb
&�KM���K4	T,$���T��SM���Y�S���	db��:#q���>��R�`�4�~��k�9x
� Q�J޼aJ2m:&0��.�x왲��F������	���9\o��l�#��O5���׾<��"	���cG����	7l���IS;
a��.�`��AVH��uN*ɛbM�@y�&�̳��4ZQ��5��oY%���M����͖̣��l������VEv�j���T�sdOof�X��9dt ��T>�5�~t�m��J���;���B�I��ޜ!�W�����_�zT��, ���%��üx
'��f�T87��E�R�+�:�w�Dp]���L�e�����P�"����X���j��H�֩��E=�Mf�XKg�|3Vp-��\q�>��5�ԑ�>�idV���1��q���(��#�@��B���IǭMP	P��\� @� -C�L�=����Q|�6>F�������lc���Q��/yV�]Џ��3lZW��J�m)�p)�tw[�C(��b�Q�-�3��ԓqO��2;���lY�j[�y#�郗x���g�}�l�p�5��yJ��jF/.GD��*Vk/T���{���[�H�<Y�I��h�zز���ʹ�p����vz�>G����щ*Ӊ�qz��t�G9i>xB�.r�hÙ�5�Ĕ�at�og��O�ٞ'���k�~��@UM�]��m�ͫl�B�T6���H���|�Ujp�sR�"��Chե�io/CR�|�e�v�
������'dv	�}`��DbX>\�����]��"�Ea�9�T*��� ��z����)x��9��;J�s?u�_�@��l�A4�">��:Vy��-��K85�^��~�Y���X�:��yVܾW[6M�����铴O%�7N��ǐ�s>u�0�]�<�oǹ��6:3�	0�T������iF���������P �Y�x�U�O[+��C>c-�]h�Z������C�	��6��6vϗW6���k7��nW4rಔ��0vk#i�w�.�y2�"�3�W��F�ciۨ���[��m���[E�Z�r�t�B;.�Db��6�tR�Y3IFe��ȁ-�����~�8���`N<��'G�w��1w7����d�ad��#W1H��N�ǽ���PcgQ�0}9'U2�h&�0݋; ��+�U��Ew:ۂ����Oy� i�ag*S�1l)��/��q�0�3����lqlB����<(�Y���8�嬮���ѭ���R�$\��	LT��o�,�[�3�Y�.��hݪ0��2C�f��T�{ay,eD�^�������v�P�'��~m��n���R�Q���@��O��lg�8{�T�=�)8�x���S�"`�4sȗ��6s;V/������:$q�%��5'��7g�Mwb��E0y�}6vn)u'gϰ��=�ϔ	�d���9�y�����yv��� ����"��7|y�ĥ�S�~�b�S�Eւ�Tq� Q��TR��n��tO�|��\�{��-C�q�s��y����D`V
񝅼�G�Zoy۩��Ŋn�Yq�φP���� ��� eF������x�In�+�M�'{�2`bs���+�A���%C�(ϱ��C�+t������i��
&?RÒ'W	N�L�G������E���m����_��}������� �e^���+
#'ߢ�t���2��{�"a�`��f �"�v��m�����W�J��O�;ivx���T@�Υ�B4�����&ɱ�_���?�߶�>?��Q�	G,{N�b �d����ɕ�L�&Ѕ��aJ炡ԏ��4�4R|�� �p83��ڜ�������A����l/�\춐��S*[�z5I�F[�7���AFҭ�E��u�M�-t�F\���wQ�N����ͯ<����*f箸o,�8X�N �x�)�K��@��y����I��`��K[�9��"�T�J��u�r�0rJ�p�flX�c�U{O*����Llm��gR�fL�O{�bOB� ��H���
~�,��W��$�C=�l1�w�v?���\qv�)���C�IH$V`.'9͎0�w���A�F����N1�J�.�t�s�7�4�J0�c�ziaan~fX�\��m\�+O�� � ȷ��?�D4�������7��j�6	w���.:�*8`�	2��|qX�c�Q��q	�����'��jn Tj��~��� ��%o^�5������
���2�l��B۩M�&ǐF�$�cC��Z��S�vt�wT*�gX�b[7���`�K�������=~K5D�̕~���$J�?=*S��en�o*t&PQ���2.��k�!O9��r�e�����I8c����x�Q���U�oƬTi�	���ω��������\�G:c�<��6��G�S�4�����o��8~��-yP���tm!u��M$��
V�Y?��u�T�Eve(e~���^"h����l$�Ef�qp�Ub�����&�9���s��P���+E	�M�>YSCՃ%-/��s�d�j5?츽wL��Ar�����;[�g������f�k�m����.`e:T��q�><7��h��4c�r�5�T�ʚd���K�bz�;���^�'��ɗ��[28T�/j1 ki*}82{����L.Cz�)"��4�ajs�+��}�8	�*,�!{]��d67I�gf�L���g�-�5���pF���g��~�UF+_���%�Oor+�Է����R���E�tO�[�-��.��,�J,r � m/��b�c8��ӨC���i��:�6`<��>��	
���k��"r�f� }��p�����Rs�Kz�v�> G`�W .�sF�8�|V�����Q���� �!W���H	�CȂ+�J_<��-�[i6#��`�"v����%�����>u��y����[��)�X�OG���]�-
��1~�W�d�m���uy�����o*CYq\YUf�����L"�Lk�}����c뜊s�qe�1�~22�!�4Zt�Iy���M{� ?��9D�"M��Nng� ��A���X�hQx���I�
�	a�[�:�g�<�]�G��r0�U�ru�����Ӄ��?ň�^R?�//�.�����-���x�:aR�$K[�D�+�U��J9K,Į�o�F��)�<�m�[W��V���Lf�:t�v�����-Z��M�0����5<��wcCSL8C�k�$�>piI���1��8x��2SD�CN�����(V�s�h�z���\��
�v�k��0�6em5���D"��#��-�R{U�8�YA\O�µ���e�K�Ȼ-_����&g�w��u�kḬN��O�¶�Ra�+e������r#���%+��NSV'�E�K��������萷�� )B@S��N��cnK�����C^��q�K����w�k4�L@.�����ğEK0��ٔ�� �X����U/�U�r��̙H�n;�9������$��j6��Z��Wi��?����]�Y6˙\�Y-����S5вdy���y �N�b(�݂|J�T#l|�`~m�.���<8�+K��DL3��E�=�B������12�:�Q�8����	�ZG�pj��2��F~�t�2�T,F�R9k�e��}��Z�QD@�28� Ek����Z#3��TB�9�F7
���Եw~���� Z�v́�@�a���_C�Hl�

��-� ��V�
AE�x��-a>�����T������=��1 4Y�n ��\s�
�!Kr���J��� 3����&��c�ΦS!!�x���X:^.����	����+��E�{	k����FQ�L mVa۶h7��O���B�n���"Fs����}��^t�%�l�HF����"%r%\�9W�K�+.���ӅHO�j�[�T��HPu:��Z-��&'�LQx��$TE�K�r��mMh�a��P�&���z�dks�¥X�`��8��9�93���!/��i�d�C��O��������v�Z�d�Y'�_���sS2}��lf��X��8G��vc��Q��t�F5��v�1��]P-)#V��%�6�O)qz�}�y��-����Vy���舞'�f��Q�X�qj.Z�6�L͋Q��rYCS~��o��N�ZSg�D�w�#��~�~:��� �M��zN(Zx�����jT���)m=k����y��2��ئ�kT��Ο$%��5о�n|-��OIcF�/�Ə��R>�����H��\��2	��m�nA5Q�����"�I�]��Q%�@s��z5���-�BiX�d佥���V<���B�pb�&u0������Ji�������Y�M��oȶ� m�ߓ%���U�#���2`���+v����Ɂ�Dӆ��a��/��.�j�
�g�=w��˖��G��Ҷ�S����c�z/�O����7+A��*hn2D����y��9�d�^�~���j�4q�Ga
�]ʓ�V4�@�������Q$҄����۠v��&\�-��kW�ƭCv^y$�O��.U'�9��s
߯�!���{�0�¾B6�t��6�'I�&�QED���O�1�&Kt<i�"�]��^g�e�Ř�j�Q�+Ͻ�$���𢢢i�H�RH�c;]����NE{NG݋
'�a�AW��:��xeZlS�;��G�.���-,W���� ��MĘ�H������!:N0o����z@��+�:��;]W̨���Y��2�pϝܗ0P�ܶ�L�j�n漭єŲb믠�K�=�;<e��������۸ä�&��d_6��g���ީ��z59�ԝA���P�۽hh��[J52�-ld6"�/�Ѫ������b0�"Fț�"Ӫ��L��b+�>)���{^N���J���ʤ{ɷ��W�R�;s����Ŀ}`I��KTE@ a��ѓ����2�v���|k�z��U�E��en����
�J߱>U��Ѧ���ªyo�rY���Yr�ټ�������CH��*Ƚ;�x�ꬋ�]*#��h2M-ϝ��`��*���l&�U-g=�$�G��6uL:7Q|j��g��v�8yh$�r"[e���i��s�w�?�^A����Ps����ex.�� |��<�q�b+�W�7qR�<|�T+�>ˮ�"jP�͊[���i�f�7{+����6C
B%,B�(��9R�M��7�K��4�� pzT�ѧ�y��E��A�!�A�*����$� q�D�ג�
��՘mj���v/�>��p需�,F�[�T|/�{k��y�:��캌 ��M)��y��ʊn�}�w+�Y>
j�[h�����\P
S�~#gv���$y��D�=�1�nhd����p��(�j��`)�/�����`�ǂY��kL�;�|���k'��0�^P�e9�D~;�0n���^�ZD�����T�'�����ED e �h�_'����}��Ay-;��Ex	Dׄ�W-���v]H"sG?�f⛬�"�}�+��b�E��h�e-	%�M���^n����E�����ѵ�)�ǙC�iZ�_����J�+���_���
V1���~���/�s���
�O���P�h	��v'H����D�nn��_YI_U1���}b�2����Q9������uؠJ����D��HW�$`�	�"d��ɓ�,JQ�7�J���M��:WG
���Y���w_�	*5�M�z�<�����f�Fv��w��;! ��h.�:S�籼��ɏ�~�5,-^a�e��Q.��H�*@���#��ڀ�q2�'�={���Zp�D�3?�ԡhٖH�5�����(��˧���w�7M��P'r�6o�{ay�\�� t9okwk�Oe[o��]���}��F!3�]��tqqcs]C*V3�}�ۯ�Q`,q�B��b5��gh	�P�=4��z� ��"�_�������U��S���wp9$I�r����1(�Gg���Ϟ�7�=�n������?0}mYsR��!���n]���<��ۚ�Wef<@DI�	c��
S�^��� .�U��ث�X�MA߁)���3��}������LV�=L6"
̪ _��Uo�Q���Z�����*s�;v�c�T�9�&�Ӏ/`A�� �'���S�u�2D��=�\\ɕ�ΊTC���g��*n����#J�!ïF���*c0��t�Meϻ����-b�� �WG���99�����`ܾ����&����X#>�_I��mA�o�ƮC`�[�#��$�^��d��P�⣪8��� +OGEH
O$u��	���U���|�½��()��~[`�_VC	��8�Y�A�g��)_��f��G.�a�.�Q���m9-?���?]!)|I���4
���ፐ۝]3�!� ~k��eV�ć�U0"�,'��7�z�Mg߬�$*1~b���10��R���m�JV�n�`��jlY�k�	*AX��^d���8z�#��KZS�%%���i�
5_�����1\j�����6N��$<�Qm��^����`�p�q@�@�!�z+`��X w��J�L�GU�|���0j��x��7�&W��ux5X��pT�݁3-��K�i�|AvF�ąՐ5��aC�;���3�� �(���)%k��r�kX����R.6a�,FN�+bi,�����@��
��6��̩���F�±�pat�^
'��<���������RT����K4]vo`�x�J����TE#��3�4i����=�H��F��n�����{�2�SGRpzP� ��q_�״�r/Wz��y�J����ӈ���F&�Y�$��Cro�,�+Z�hg9�}�STX�6J��a��0���A��N�3��l�u�����m�T9C'p���H�g���Jd�
l���7�ÓHEz�`��[���Ҁ`�Ir��-���x�RAy�E����߷�O���'L�a��CCi!,y`0Xҗ:27I=�Um��A�q�\����T�J,���7Z�Q�)V�V����~��?Uo�Y���N!��էZ6��MU��;���$Fwx�J/���Ĩl�l^|ӈg�2D�6��LǗ>�{,�2'��[Ǽ$�����닽Iy���b������o���}��4mk����=r�=z�� lSd"��5Q��,Pq%5����gO��	����M�9u9J�G|ֽ�������O�E*i�ό�
w�Pt1����(d>|���]�_-�x��!M4���N�I\`���p뻉�Ͼb}�A�x(0�
>p��]2B�1Hm��f��x����	Nڌ����Ǐ=A�����ph}v	�>h?*�, ���:�A"!��S�-���H�G#�&!����f%-��1��}��(F\�Ŝ1Z7���X@m}��"��v���nz������wU]&\0
��l|&S=����hn?Q�6i��1:>t"�\����fҕ�˰n��A�$��n[|Ҕ7��ɉ@]��LJ�8����/��`^���tY���х��R�wjC|�ts��^1X��'�0�lTaa�g�m6�����Ӏ��t�ީ>0 ��*�Q�@N��M�1.<Y��C	���g<�c�t��U���Ŀ�y-�l��sz\�똖7F[�Z�
�P;h��Ѿ�J��0��N~�)'�oY���c��O`_Sh��t�N��z�Q����M���ON��b�}��q�ZY#��x�8u��|ؗ��C�(���ʦ糲�i3����>�K8P����&l������~��b٨����ŦμzP�Y1%tD�������B!ʷ��M!���� Yd��g��x�u����,m
��)Jt�� y>o,�(�-6X�ƿl,O�-�"�Ȼ��$�����c:aB����w�74'��G$��:�S��U���2�Qx���
W]܌��E�f�;�j�ϕ4(����jI�b#'�Ӡ�_O�9M<������hRKݚʅh���ƾ�v	j�[�sh�V�>C�L1٭<��g���a	���*J�VniJ�gxA�T�~�yv�Vt��7��&��� ���N��p�d.���ͤ꿻h}PC U�[߬��� ��d��Ju�V=�yz��CmfC�P+6�^ӏA~�n�3��n�������y@пK�-�s������d�fa�hcږK��ғ�|�d�v��yi�Z5�i����C%���8�P8�lJla����Hy�.����q�*Z�o�%OX~ԋN�jٰ���&����p�����(^���m��Hɾ�$YLrA�gܴ�4��F\�b�������@"=
�^v���A�1�|ƿ�pIT�U���y=�3�Ω���+Z�s0�] �zॗ���6�K�:7�<OD^.߯0a�Q�S'*�E1�Tn�<Y�@dIh�0��?�Lct�r��!1�ۜ�ݪP=֑���Vr�Y������}�������$����<h~�Mt������\<=�݁V?%��?<�ֆ"̥�A� ���
��C���<��I�Z���gfLJ��w�j���:A_ Ϊ_@��$�Ie4�ցRW�;pg����5+�(��ѿ�=�n=Wf��M�"�z��Au.NzoJ�����Cmp���r0�}�0��o7A�R�P���s6��	QG��߬z�f��7�㚭�y���/'s�85�V9.א�<B=B�0p`�������hj�F�֏����>���鴼�U���K��fpog�������|����NNip��T?��?��'����C,#��ֱlh:�c~h�[1Mm�jl67����cui��br�2���{��w	�І��Es�)s�n,�?�ӏs�fO�����y�6C��G`�,Î6p�x�A~?�ZX2�g�Ǜ
)��ͭ�E�·�۞���
����4�j��{�.�����I��ٺ
���65�j&��'��'�,o��
�Q?���U9��buL�?ٱy\+75j��MB7~���b���c�G�J�h�g`NJ.r]�7_�HPy^�~j�������ҥ���s��,�� `L��n��L��ۅ�!濒��H��޼�	R@��Z/{�6oO��W� U���l��^)}�sQ��I�+�O�Byy�_���.�L�L&�}�U)��$
}o�U�*�9A�/	& �X�u�(��uI�E����v�ͦ�T5'����F�Jz���kR�|��_DY��
�`"�I�QNv�kD7���{\`�(�8��*�b;c3��"B�R��$���P���u4V�d���d�,r����q���Xԩ��È��L��=�[�	�r���P�ȅ�A^Lj��I��<�����ϯ�\|�:��!��a6����X!f4a��	&�?J�6�e0�,�J�����Uҵ<�"�t��S��7ɺF�
S��.O�Sm���s���>�ӻ뀞�b?�<��5�0�wA3��2�iK0��:i�X���+ӭ3��I�oX=� �����2���%��?5�Ej�&u[���M]p�E�s�V�O�Q2 OX��x�j�	��*_N���31R+�)��F��qo�a$��X�,v�i���s?��|��1)w��ec_'�}�����p�%^��f�$�\��)�f�� ��\3��]Q��G+h9��;g��q���#
7��qX1+-���J�n�W���f=�:��c|��$Lg��]FŞό����gV���{�B*;89-^`r0��lr��m�eAB	~����?Lw��@�F�.��}{X3���i�"�,�X�kJ���0l�޻��o�)�6�4���_�(�u�&���#��*�p+�ޱ]_M�~��vE��ݮ��%���GIͯ�(}�+Cj��-�R�+O��\X�	�O���6�R��o3λ�[���8=	���ԯ6���3�>��`n���o��L� A9�x�F����֠6� 촱�o*d8[(���j����r��'D3X��/���9Js�T�NP��������I�C�M���գ�e�Ô�/��8_��o�K�Y2�z72[�!z:�D��ƥQ	��CB]Yn�Z����[�WX3���Z��`!�ה~�Ch���������g#�9t�l��ެ�5+�H��X���`F����FMB|H{sD���������ϲ%�@���z��&�8����΁F�hI���Z���Dp	�i���S������q��1@���[���EE3zZ�z�]�%�B����ǫ��1���8a��wT�H���L��/�٭7���B���%��)�c�փ���H+���7!�8v:�^ �4�ɳ�Q�?@ ��W�˙l���{!	�ܡ�͔"@������l�����76��l�dtM8���7�[�U���S���+��:3wP^ݖ�y$�y~O��� ��;1�M��J��]���--�ԉ�N
�6��TJ�Mb��d6�U��.���&5+�%����σM�c��$e%"�p���zJ#e&� �F�P+
9����W� �驌m  ����7+wZ�����t����F���ׯ�~B�X�hڡ�I�훂k<�e��c�(9Ɗ����N��b
�#wN��B��о��ʔ�s�b��pk��¼@X��l����F�$��B��.�O���&ZHe	͖u���?J8Hf0������Ü���
0 ��\h� ��o\����{�����Q�JS�Bb�'��R���zF�Z5��cl����+J�*Qk��2A*D��-�1�*1I���n�R)���F�F+�B���\۶���?[���ȩ�� ����Q�Fٍ΍�j�TDD5M�ſ��g���ϊ7��E8��T�V�$�S*���q�n�>l��րf�ӄ���vP����R���)�0��b$��@s�iS�]�/�I��`��/\'nѰ�I�`�U1U@93�4��=w_9�״�W˓\�dk�3��9����j������fB�� L�Q��:|�^��qA��K\ڝ� L� Qc~\g�~�m�(>�r)��-��B	���vꚖTO4�
�������\o�h���p��ɔ���|�����������
3���v\�k��B��,�M==��4V�
ewF����4\�CA̍��ݿ'��s7�SS��i o4J��Q�y���>I�z��ſ��{S�|�ʹgq���+��s� �3��X:0?��N�tx���4�Q�@��Bc/x&4_3G���5�0�H�{�͕#�Rٍ��*4��=�s�{W6OK�+gs��|�l�}B�e�iό�*x=W~_�@:�D������J���ў�Kʩe�����#�y-jB�����3%d�'%PP�`��/�6r����+��~w!>X���QMҷ��w6��eS
c=�C�)k�H�p���
�A�Z�QU`q����0&9�h�3۫y��uZב��Wp�7}Eփ���)zW�Ⱥs�e˹�f�s���XL�<G�����{���(*�V�h�gt4��95�G&�L��Ҵm��X��P��e���:K����@�{��/�t!�Su��u��Psʰ���#=�ss苣���p �;��V��0�Mn�P8���	f"����ؐ8�R慳@{��8%����m0�D�H`"�@7� �=�����ý�.�ԥ?�ӊ���	N$���D��6��02�9e�>�FA�M�}��x��\��.�L>���A�q�ʘy��~IC�w���{ma�8���Q	�͇s��Ԟ���i;�)�s���/C�a����Q��㞠-c�!���G��yA�	��͙V���aMҧ�����93Du$;���s�u�+��0�Juqo�åv�J�W?�2A�[>��=��AR���M�E�ŋ)�lՌ�.;ˬ�`l=��Z�В���F�g��
y1:4�����u��i��"��,P�ᴞ3��2&���"u�iH���Nc���J���UJ���*[T&�������^�b�!��ͯs4.X%����ʌ0�Z�A��9s�۵�~(n����H�����zHp<`Z/����!�;(l���+b\�� �,M��Mx?�F�Pk�t]hЉ{s�O���̗QM�\�FC C�.g9�����+�7]�����w����1�f�Gp�#�Xd���yxɟ��#�c
j�H�u�3�-�&V�#����_�-Z��9����GYG�����|㝸�w���)�(���p1�+q}�*I�|���qő,B�Ӗ>��q��:�N�2Q'��CY��[��^v���5�ݭ1��|q�%ז�����;H�m�	�˴��0�-�������U��)�-xr+�+��6��=2�byU�([&A"V�����TQ+���R�CY�:Ԇ��ל!������(��(L�5mn!��+r��_�|��[���;�������P����:(x�Ė�S��U&�S�����'ٙz�IFkwk���Xj����}!�g��x vG��0�h�fص0 5�!����EW�n%vC�u#�?e�-�Cn	��
�ـ�>��	�>��{UQp��RD�{�h�y ߙ~$�V_P���[�)�bi��\����M��z�pgZuGj�e�.Fh��� ���!�����A�GtT�<��3rE�8
��z�O"��]���۵��ۢ�L�(N%���(#N#+Ҳw�sֈT�#�F���xof�&�β�i���x���-]�6� �D�r���Ⴅ��0#�f�zЩ�W��aF��K��{p5��ǳ�j�ӈ:I��� �\�;�0�D�[��F��@�b�`��X����:�q��zL��o=O�A\ٲ�/��Evc�4>�=Ȃ[<(RW�@�}U�w?�|>��r����5]j�{'���.@�&F0��3���4u���A�����f�n2Y�zb�|Ɣd�[�%�'S��b�$!�+���>A���1��?tk!� z>*8��f#`,�����$��r�vr8��GD���>H�� w�A�8����V@�$�)�ޙ�ve��1ď<��T�ڦ$7�Y��J�g�N9�$��d���}���Ro|P��.7�=L0jxH!P��0_��?�YF�غ�U��jy���m��pHg>AL�V���0�= ��h�HY��#�QT�O�_��� �}B�	{� ?�8�������*��R�� e%!E�i�ΕSgn��v�_���`�F�r�V�%|����$��}�g��m�e�,���ŽGT���By����z��Lb �?f�������j��*I���b�lƉ�?����?���L�#�"�RD�&���yi�S��*��ձ?kUS@Qm��)���2�L��Tp�&cE�y�+�
������{H�M��6�pΛ����M�[����1�eec�U/�a�4�I�*�͵�����/�wod���(�]�����]�{Bу_ر3�݌P�����D�#�Ԋl��˾T��x��eb˘�����6|�*� �b~��U��%B��<�c�$h��̗���gB�jL2���&���0S��R*Gt�B2������+2س|��Dڿҿ�c��~��}L�"��RW���{p/���J*��<D!3�a�b�=a�@a+����;ą8;��e�x�G.p/�ć����
h���CM�l��_�����y����V4���%T����J}�t�,�ܵ�<�#����b �Ïqe��'�ɕ4��E��y�1��*���y(�ڲc���E�f�7�[P
����Hݚ����Y)֎�g�`��I��ߡs(��k��� ��*V�^L4�=l)R6����S�#�^��|�'�v��=\l���\�Eu;�kA�� �h����m���,G���Ͻ���yA����Ur�Pr�9Q=���-/1��>}�Mc,~W���G߬p���s�c��s�L),�e3���^�堨�֦%�6���y��^����Kj�sG�Ϗtd^;��Le����g�rk��R��eA��o�.$\��\�͐�T��П�-S*�����>V�a�����$��T���h��2S|�!SD+n;�+X����N�M
l����ڽ&Jr�4nx��e�]KK�A���	�c�
�p����{X3��qµM�x����{dl�x�����l˾�C[ޠ	�ߓz�^r�"��8�����DOR��M�ٽr�F����~]�
u~|���Q�@^w���]&,D���l�v{��U���|�*��vHR2���/�"�zuQa#��Se��u=����9,��n�����;��+����&�`I]�_�^B�ލ]�C:��Z��_
�M���Hp�mzF캬K|<�m�1�r�kLTh8�,-�<�r;g�A'�P�����Op�j
޴�U����+�cl.!��3̃��t˳|�/tl}h/��!�0��o�(�q�8֥M������>�<�k�_�?�=Ϫ���X�c�a�F�k����<�X�؝�� T�o6jH*�ޖ��eL'f�k�f�d@��Y,g����d��M��֙����}�1�\ۖ�h�%�4�T�D�V�tQ�67��r4���U8轑�r(bnE�������2�c6�+I5�K�5-*A���ZҺ�4��΅E�+��S���.�w�[JE��� ��%Oz�`�E]1�o���M�A���%f�&b�����
��^&��˝�+���z����[�3Pk)z6}�E���ᢩ� �G{ot06��6��~4V�b�Ԣ-Yk��Ϝ�+[V{�+�r�w������ l- �^�l�#���:�.�����S���`^>����S��ID�f~x�;��%��\�:�c��=�&�(βN=u�؊o����8��<%
ؠT��U�;�S�b;�~B׏cu���ܞ���~81����Pȏ��%��r��r W��<�@�Ö�P8���[�)�=�E��Q9����O�|n(I����/���"`;@�rK2�&�[��f<.����K���'�����M?���}�����z�M�K�:�@�d�U�w��g�c��8���&]���?,J"����G>��l����S>��Le����*�1����Eŉ�׫o��rm��Kl%�$���Z�$�Z(�šYMk��&���Q���N�O~��`�v��+q\����dY��|��L�\����
��e��Wu�C�Hy�إ���t��C3�&�GX^�v�*P�%���Δs�#8d��}B�=�c�7�S#��+>����%d�����J_;�l�X�\&T�6��h N�Ag��� �zG�S�.5t�\W�S�{?0�x;�j�b�2�86jG=q�����>y�zZd�'���3��g���KG��d�p�7&������U���i��2u����W�$Q>Urq�@�&��ѹ}�X0'�9�5|3W�Y��o+����Pì%�����0R��N�tzȻf���*z�NP2����!0hg�`'0{@��k�R�I�z�%?ia"�ȹ7�?�Iˑx\��P�KYC���ӓn�T��Jέ'��b(k��D-Wٻ-��=&�
��F�g	���|�/F/ �Oz�m��j��x*�����?5�#RÄ�-��6O����t�E���m�6�״V�K�w���w��ġd^�rg12��Nlӆ�-i�v�~zf����UdIM~�`�J8�����\�1}��X�	�����`�Y�� W�U�����%פP#uv|v3�S��<=���V��o�L�P��8m�O���=�����oZ��:�i�@�򚸹��=>!8��\�����~ $��<���O�'��O�qy*�-���H]�w�&�If�\�u&�e}��h@�x�Y�Y��{����>�n�\��:��	���6��o^Һ��*a�៌w���^���ʑ	������-� �7�9�&b���yv���U��s�/�x�&����;���A��s�����erϯ��&y�
�a�6�%�7�z�d�W��n��B֗�ͧ.��Pl%��~�"��VFwp#|��\^����$��1tA��"�
����ÏO0�����A����3Q	�$/�gӨzc��2,4�^���@�)���d���W�g��_�|�������|Q
�#J��r���:9�_�~��	�gB��nRY�
#z�E�wTSi��F��P���Q�x�w�G��M�A�Q{���!S�4����[xvXc>������]%z��p/�ៅ���9|�\rl?��������*PASek�L�F���-@W ���m�p>^����J�HbM�`�o��I�h���9�+������4���Lކ!%�$Y�P_2�)4��xP|J���XGzK�����59Y�0�m�
X-�c�C:�2)�{Cm!'��f�e��+Ԣ���Wg��e|8������DG�p�]=����X.Hz��~��4��9z
97�R�Eq?q\��V�����z��b��TnqL������%��L�[�-����ƺ����8�*zB��^��G	�u����������gz�Xd<����^D2I�䜴��1n�W	+J�@	��\tZg��dc�UĊdf_f(�ߤ�b(+"�<�܌M�R�~�.���t�>p;B�a��c�@W/���l#a�0u����̋�V�]�zg�{9��]��G�6[ `��3gԴn5���<Ù��p���h�c譻c>=��	�9��<`<Ѫ�:PŦ�˄"a׈�0ε(Q=�c�Ԓ��P�]���4��~�'���P�>=�K�)� �[xk=�k�1jT Ǭ��?%��Z���jI��Eۨ*4�e�кz������7�8��)߀p�'~��>�(�Vu7�Gw��u8FjRy�	/�Ɍ�A��Wd�-�����\�2��߉���:��@��ɥ&��bu����̕��R�3Y�D��'K��Lk��3kL�1�W.���Zm���8������G�ٿ�&�Ixia�6pV�埠�O-�fNFL=�km'�����')g��'Fa��MCڵ���S�<��*JZn
$_�c6/��,!��t��J������b��H�X#���w�zZ��iѸ�B�B�0T�*��}�~�}��H�"=��s��_�۶��Ww�?���\�W�y.��c�|�����*���.Y���3�!��7kU���ɥ=��B�}&��ް;��2����1L�tޅ��y�@"�����V����ǵ	L�S��Lq����^�!�v��~ٵd�s���ɪ�/����k/�{�V���up��,:�m!��x��r��� <	�u˽��p�zb���Eb�ig2��b����h� %��I�-�9*�9�1�i7̬�3��jA��#�ߴ��{fC�Ct��0�i�@0C��#e�n`g�#x��P��S%����l��aˍ5���1�!&�w���f�rmݴ�U��^�ݾ����o�:�Fk���}�8�%���_5��/�Գ*ҍ�!&@���+R�ֆ�'�O����@�� $Gx/2&����c|Eu�: ��BM��Z�O�`*~z�갬P��2ѵ���ﲦ�!jY@�wt�+G.x-�鶣�o� W��p�ٯ��0^!��8� yZd�Zt/�ZV�\dV��f���Xz�(�:�����<�$����?�{H�7K��m�ZiX�r��4���8�����|� \�yʿ�ٶ��B|r�|d́�=|V��eajίg��,S|����E'���r]�K���t�,�/W&&ޯ4j>5l�<��[�hk�P��(6l/b8 �8�Ƽ�!C��ϾB�:u:���v��z,��`�s�p�_��e���F�팛���X�>�2Ц;�C�]����-�Ii�(��/���Em��c�GN �P�{��ٚ�)x�z�9���D�|�4��ꬢ�n7�
�qz^0�r�d�Ž N������r��2�(�Y��տ*s�}��*,�@�,���.����r����84dJ��{xs5
�՞l��~�ei�VA�k[-�J��|�CE~A���Z�N�ihu%ڑl!�G\ n�hX��#��Ǟ�s{˅�O����/+m��x���ilpI�?��ӫK��c>F$���E⥪��ƗaB,z��`?��� t���~��_����ʂ]PQc���$X[[u�s�|ޯ��FY��]$��ک652��ܜY������HSy��<�X,�A�����?8<(��[�hH��ԋ���!���=�f	@�I�����MW�yyg�ۑ�'�z�@���Q�
t�1U���%�Q�+jB�sD���c�t"���	�KV~
/���Ie�m>��"_X\�)f���{_��ﾠq���p��4�V��e�e+�1(�y\�1��QOz~�vh*�t��cU�l	Y��������<��z�M����y�[[1Z��x֣�U7%u�����b/'�x%�>�����|b�IED:��&:}���XC�4Rhqv���Kb��'tG&yN�J�)z�<��g�*��Ox�#��Ԉ��u����P�5T�;�/�K���)X�C��4
ށn^��x74y�JB�\��˔�D�������F|F��ب���H�`���֘qP_�T�%N�-�-�67dA���-m7m����I���Y�d��c�����\��Dc2,Ѫq�_���K��*'��si|��&���L�,GTP�k5)nN� �ծ%�|�;���^Q�4?/9���!�Z��,G玖b�]�]��ˊ+N6�~�r�j�-o�%gu��)5�~���#��&�L����h.sӬ��8��#�eې������QN�It��r�+-M������>�\>�BMz�y�����'_扜���?�К�.d�Б������`����M6�K=q��z���%",�{N]�n���ՄW�����w���'#�0n�����mI}c���I�O�#9�a��Pc�S���,X��q��ۈ7(�,�.�ŵ�c�)��X�3�Y(���Jf<з� �O�b��^v4�\"��]Ǳ��O���`0�h��ǖj��ٞ>»E�M�O����d�} 7,�ݗ�����Ac�Ip�/��J\W���^���fV�@�vZG7�r����M������S4}�A�K'8��@x��� l	��C�i,HZ�֎�MT����fK�[�R/���&�Wt7A�(�i�A�����˯dPV#rS�_F����oY+��p0���Z�.ĀӲ��2iy �K�p�XwS;�&ƫ��oT��:���5�ͭI�R�
ιԗqb�B������,4Ҭ�WZ\��=wt�;��N��q�
��krc����~t��7o��*�_/�C��+��H��t�5�E����_C8��e��8���B$CsSim��K�W~R��_�ƗS;Є�
N�I�>���#��91�)���c�8>��Jw����Y"^����%�lyG�-�.����8�8L[������qi��Zt��u���y��Iz{�ž
�'O���Y�C$�ۋ �u�i��V��q���֜�߲�#R V,@H�dd���yy� �K���e�8W5��EX��_ߛ��8*��qjs%}�I�,��ӫ�c����UӪ�,5N1�[��{��&%B��3M�@H���n��N����f�,��vN@4Nn���H��H�S�}�?�N� �?s��(��g�5��͙=����S|�Q-���1�E����B��ش���v=+Q��]�v�g�٠ֺ6�҄5(A��ex�`)�~K`ӯ�b�#��%H�������7k&�S�g&F����G^~cR�~��W�2֔gA��q�O2H��@\�%		�O�r*g������˦���M����TPC��eC���t����Յ�N!h�5���2���z#�V����kN�ً�3�;x_�:�}?l�57B^�����Oi<���v~(cQ�PQ1���1��cvԘoT$�`M�)6NZj��d�$4s|g�t��1D��'�p=��n�	��!�� Q׿q��53���M�8C%��0��򁶷O�%�1��6؇��D��D�ȴ�����1�0ָt�)�cXX�k��s���5�D'�L�\�FHV�J�`�@\̇�Nnbt�SV?"�u�|���Q�UX�D]1�
��=_�1��)��.�fD_$��Q,�sq>��(&iAG�I��^9}��QZ&�1���˕�b��K^\�)B{�n$��~�8���s[���hK8���_�:��:�UϹ}Y�J��8#1����v榊���V��e��/i�6��3�&'��=�y���9P�Wm^���а,�ip���g����9���w:��%^.�l>6�k�`��֟<��Β��z�V9�C[�[rwM��zIg��Դwb`� ���6���M���ܹ��=��}��G���ZT95B�fLd	/EZ����t�j�_x��h����C�V,"��y��z�D�jYք W��/�+�k�I�b�a�}ҋ��4me���$Mǯ�堶�ԧ}��Ƞ���j����O?��2�-G����o_|��Ar��;�
���}�>�B�� ��Lf��ϛ��u-rӸju2Z��Q��`43k��'�
*�I~D�i"��i��B�R_Q�1��R�c!�j��ǝ���dg,���_ꡓ� %Zh�ӣBwb,�[�yǂ
y	,y�����^UJŹ{���p��O���^P�5�)�h��%�w��cD��ȣ_9N���b\k��^'r�F{N�%�{��$���'��Q��4q��V/���|���%Z~4�F��-� 4&#f���X�W��Or�� n働=-?|�pH���/m�s��#|��k�.�m���Q�!��¾&�w. d&��V����d�p����-a#e��rI�V����8A��t�7�Yh��O�MA�*�1��:��Έ&��@���d��Y`ב�\JY����(2�sK��W
�J4D�v�U����n����H���I�Y:S=�����t�gu\J6E�`h.4fj��3$�E�P�`�p�t���g�ժ6�=$tXD���J���|��nh�YC�cQW�k�Jտ�'��ʮٍ��Ǩ �}���X���5Fr��ӊїL�L�!ev܅Q $P��sA|~�غ�4�*ݘa躭���(G������j<	�ʂИ��17�¬}�#>*q�Bۍ�5���X�X�U^��-�{��w1&�,QF�-{���T.��mw�����:����(�a?�K�����#��k�0㍏���AG��!����2<ţ�j�<�b�a<��_w������5<���a���S��7�c[+��a�ـ����dЅ~A܅7p%6E�H�7��'�3�?_P-��ʅ��&�Sô�`=�I�5�b�DQ�� ��rمV����敓4� �Ɇ�o,_`�<���E����?�-��)����Z|�`��S��N�I��ϵ�i�"�L�� ���(t�KŜ�8>D��I��o\x�������?��H�ʥm]8���8+�iu��h�_�C�G~��_]W_n�����s~wJ���W�>����Xό���W�H����h��D>)\���
���4���lHvhkY̕ӵ�d�����eF��{�\�Ot���B�����<�&���P,T�����M���^����Y���θ����*�X�SV���Y!�? (�&�L���qC���~~� c� -|�ͫ,��D�/�[W�d'!��]@Ƴtί.����>{�>tPӺ��#����lTG�>a�_�h�C	)Q���"��
@����e��t~%�3l(Ae��,�ڝј��b���N���A����y({+����Lr��h2t�$3�H�ۜQ7`����/�*,pm��6]hT!Z:����[�rR��5�&�CG~vQF9��ԅbI�����j?��:�5_���QJ�H�vK��~��{S�I(�n4�+��aU�<�ӭ�RU���#FH��jɆD�<cu[s��2ź,�\�}/)d��W�옑	��6?�.I"�ĵI�:b +���\;ly����hr�K�/9]$-�a��(�	����Y�<|Dٸ�I���5���7� �9�(����觟Q$m/͊_��1u��	v��jU����՞+(y������|Ђ� �)���*;���
��oЁ���(S�'p!
�-q�X�c�\,���P� vg������7E��h"�ĠI�Hș�w�*��A6*^����4���"�*��m��ت�> ~ .��&�P�<�Zk�x`-oGҜ���0���>�
�/vM�s�«��R�7�(�����Y��O(Ex����I��NH�PlsG��� 2hm�m�Il�����?��՘�� ��$��=�9,\3H��j팟g*��Њ��;8��a���oc=al�]��|a~%���&a1�7aI��2�`����־��E�F�/�N;0�P���\*@�'*#iQ4�'��6~����',�����Y�d�,���=����oY�՗��}1L���N��s�J7s}-������v�S����
}����n{�"�0�6�qI�;C�ƀ/Y�Vi�p��a|A�/5ջ��F�`c�Jy��m��sJ̢Z��GE�6j�k��׆����ԾӱBX`�6��/3������	��#���]w<_H�z��(�>�
'�:-����S�p.]%h�]��L�>oH�+=A��Q7I��1�O��D_���p�h5t��z]?y������e-�Hv⮽4���Pܲ�� z������E�zW�g���ϭ_S�z�<�3�Mf�&���(�)�}��a�^a�x��QG��`�G��KR:���Z<����C>��0��W�U�Pp���^�m�)ܪe�^���GDQ�c��Js3;=XkЧ�4R��w*DNiD�x�(�L���h:3�+��jH�|�����	����r5.}�k��������v����W�W-S�-,�6	��>
� ۍ"Ox���#ݻ<䣃Ũ8/���J���m 9n[��`C�VZ��7Ƴɹ×1J7%�w��@�������P�/ڃ��g����ƍ�Fh2�_��n;�P�D=FZ�!�D�r��P[����b Ρ�5���6������J2~I����}��IM��t���9����PK���u���R�U�=�ւgr��?K��!v���'Ay�0�qB�UWҪ����\��letR��f��|�J-�,ށ���e*��$��/�n�<�^�|vU
B��5�:i�x��&!*iI���Ʊa���D�RG�Q�:��_�����2��6D�,I�k0��:���z)%��sU�_����g쿑�=�K>k�F�5v���J#p鷉ba�B�����ia�&��2r@���|5!>��� ��sz�)��s��8�{5�(�H��C4�M�a�SmP/�&��ږ��\V��(0��HU���q�*04�/Ow�np�TL��V�����ߋb��3z�n�wή�(�(�(j���l�Yd���d0�t�� h����Z�>�ϪE^��U�X���?�9���[
����nwX���ٍ�7.�]��ke9�e�q��[	����a)SE��ڌ"�p���ϕD�����R���h!Z��#^,�8�9�L���i�3G��c`�􂚰��-�0����ҭD7X$�����MWp~� Po@�2@?�f*�G�	��~���E��j�7�jj+Wf��%�Ԝ���;1�t���9"���t�'�_��{��\��u���BD�R/<��T���=�����ˡ#�"�p�l�O��ڂ�E5z�1MY��A����ڧU��у���&�f�<�n�R��Jj5���T�h)���Ǎ(���i�־���\�s��X�{"C�c�Gޮ�S���NO�i���r��M����CjXͦ�oS��Xj@@��Ş"R�=.ƔĿZ����м����=�<ID{�u���}ϔ˓2�XNE�ϔ6����	n��$������H����6�Agw,s��b�x�y�+�N��|�׌����ɘl�4��y�������]JɅ-��P�!Yf�|�On;��**Х����9����ݴU敖�5j�Q2����@B����&��9�#�%@o"��ʄ�P��l�h%�!�� ���&P=�8>�>�ׇȜp~x����e�1�6O�[f�%q�t����@���ϴS?�;�&9h�w�ͅ���bl�m@��pHc��AZm��`g�$9XG���a�ϊT`~�QW��y�S(j�2�H�7��+�ԕ�S�������du|eb1�[��^�g��^�W�(�i����r��[~tK��_�:t�P��Gy���
Bua�n�z�P��/ �G+:i�5��K
�FH�~�<��/:�1WU���n]&�����x\V�z	~�c��z(r�L�3��i�`ﱁ�*�%���F��i���K,i<�����©Ե<�7Os�I}\ĺ>�S�t*���$-.�G�V���L�� �"�E?�ߦ][Ƨ��ϖ���bҌ|V"��/��|�y�|�+�8=���w��)���V�D/+�=�,��e#�7\%٬q�n@%��G�i�y�7�귢s���@}����Ϙ���W���.��wC�u9P����𨞢ch���I��Y$�d����kT\�#}a0Ge�_���Lr�Y{e��#�KV���bŽ"��k���=���k��f)T�?|�&d�߆|ަ� �#n��#��`�{�6A,`>�Ja���"��ƪ�Y��Eg=�5A����u�g�Ʉ����������MP_o͕�8x���mg�N���߂ �7@�1^SDUG>�:E�ZH��g�8��or$�2Y1��Փ�'�K=�go��2%�J�־o�G�L_%�R��	�����}�}x- _I��%�������*S%��V�M.�$�	+�QZ,V�p4���D-J}ؼ�N�S=���G�J��uaЕ(K�w˳D�IH4��<���f��Á�w��Q��:k��Od��۠
�u�����Լ��c�*�/2�#{W��sa'R3?��}H��b��������>�S�r����|~�y��H�2�o�B������� �0�A�a�E7���^D= Ɔ�#�F)T�y�[�
j�F)Z-O^��L��9oHj�>�t�`L����T��_Y��u=�:JLh��Y��M�mOm;4M��VH_��i<��X�̌�G�������y�	.@�;����{������e�̷Z�h#�.N(c���
Xuv?�Y�/����F�?̃��� ��k�m�8����b+0S!+�]媍S����L��2Ϻ��g��>��d�5���0��k�»��*�vLeܚ��E`��:�#H�����ы�D{ˆ��/���P�_�� GO
���$�?�;�m��z�1��_e�R���$� �_��ߔ�h������80������Bh�ZР��F�[��C��?P	@�P�<��{��a��E������H���P^�?�2�X��!n�l��K'�dߵ�ʥ�w6��T�n�K>��j���8�5=rK����f!�mK�J�A}����Q�R����4^%V����[����4'�'��6o�dlՒ��@����$G{n�,�!���/%Y�N#�nW��&Ú1V����#�C�R���.��Ǿ�RHY_����7�81�M����������ķ�������+@Ҙ�_�<A>�"���Z�mV��ty�׀+;�l�
�,�ԟ�I����-���gLP>k� �CM(��$jgu@��g�d�yEO�"�N�v�������j�Vh ����`��}��|x��}��4SÁ�@6qq�F�6����� �c�a�U��F�?2�N�1$V�uS��<�$��x���!�Lp�;IN�46�4�������v�c�t#�|c񅣩�n�eIN��_��0!LQ0ݩU�ÃD
�*j��x��\L�Ȩr�PЃ��Gf34�_��J�jg�4��.���l�}���jR�����z3J����*kB�"ť;6��	��'�s�L�g�L��١y�u��o�T��ů�Mu[9�u9��.@�s(X�z1����t�'\���nd���RE;�U�o�FJt]�%�^]O+O	������¯�Gt�0A��Z�+�|�ޯ�W����KqU���QL*�nr֯	�s��̳�4�qx���)�~��	Г5P�m�V�
tE�z�sj�?W���nu��|Y VQ�\��)���n�RZ�;6N��]]��L����¥���.u��������Q�Xt1�F�_oH�-d&���.X��x��lWV%M0��)�Ix���4��\�0�n�5C�<�I��,Vr�KϏU�$NUoF�w��ۉ����íʍ��E���uPN���K� 3��5owD�RAa�Bk�������C�?��8b:�8���|�FV�ӺMS�X����&v��ֶ7�%� <�C� ]�����,!�ѹA�UA���% n����2�ݵ뗚И>���o��#�,_� Y�Zn<�G�����,�p1�H���4؎��@��
K��-�1��C{`c��Q<fO��kp=�7��J��,�bb�l�'�G]]���p�C4ksa�n�*�����5�}���t�/�	4Z�]+�<=t�F�p(e[�#�G�	���3v�	���3U���%</��^+���LB;w�Q�uc��.t�|��ƥ �B��ˀ�_nf���i�ٖP����E����f>���l&f���eo�y�@#�� �r��M�ì��K���hd�O��Zx�fn���nChӱ�	ۄ7~�8�9ǓY����S��]�YK�Zl�e�DG#G��aB\�"u<f^��}*�#N��9�Nۗ����b�W�-�BP4.��p�?����U�5���W9�f0��1(yK�~|�G!fo)|�$���V��_ԛ/��`�����@!���ST�����Za�/3�YQs1p����f}i{Ot.���+ί�p�x
C� ��g��yY�z���{��TmޥP������֤�����{v��}�f�������*Q��!���/��áq�p�C�쿥b�v�/$h�b�?�h���8�8娴�%h9�cD��}Z{�������+k��Mt�z9t�Ǐ�����"��\��g��ʮ.�I6����Ҏ� Y`���zE��C��D�]�["������[�ד���e3���	�׵�E�g`#J[�i���,T}�%���*�S��#�|XT{��0���
a�^�e@��/-Z��ݹX��D_q�ʳ@�6	:#�`!�@u���k^�v|Q����>�?�`�mJ_���V�C+Z�1��o;��x8N��T��`�+'�#.Ѳ�4��ƞ��_��'O˾t��'ڻKʙ���&ײv\����~
�(�,.a�]�@t脎
����$B�^�^���L���O�+�sG��ʫ����%�.;�L8�vk��~>Qb�`���܁�mi����2)	mw�ι�J�x�xSF{=��1'J8��Z�(�,g}�h5�)f�֛,Cq��'��g��V��o1!��WÖ��ޕR�.�t��Z2#��w�Ǎ=¯������2X������Qr�_����n�y7u<i������<��oJ��s	8��n�_�cc!�������l�j��w� -�!$��)SY黈�:g	y��p�8�X����J%�l+~Lz�ݹ��>�Ģ����Ļ	I���L��gqL#9dŭR����V��ԩ%�j=y�j� kk)�!��I`���u����i(L�I���[��^a3�֘��9�5=��A��W&�����o�	�X5���^�f�7�d�ഏš=�c0��,bõ��u	<�j���P�Z��K����!��Z���9�)��V�C�z�1����_i����?{FӶ*<9�1��Ӣ��K�T�`��+l����g�PS��7�D�2�A5��9�N���PL
ĭX�Æ�h���S��En�%^Ϥ���M�MT�Ҍ��ݒ`̦�\�����X"�&dT����>��IA�b�Y��r��TY�;�4�KlzāivZ��r쒦	�� �:U�C��g*�>�	����G��a��>a|א�/r��)�Sg�{W���btA���XK�0�|D��1��b��dQ��eS,C�W��7��u�8����Z�C�4\�_���P\��_l�����{p��̪TϮ]������^㵩���Q��~�F(�l�8Ew��vx�j�>���(��6jRҢiO�[W��T1�|s�9<>m�°�
Z��Dr-
�ś��
:.X8pR��p!R�4�;
�`;�D�����-�m3�H [��Ƞ䏣��Ѣ�����<��XA��M.�Khf�m_^�	�΂6����Y�18�rO<�p>�R�-�;^����Ԉ�Z����������b{��;/�sH���+�ܶRsj��}SR��S�,x/YO����% �n-j	\/��*s����6N,�*����������%��A{<2��!�G#��QhO�0��A��h>ʴ��3�St��;I��x�]��*�Z�۞�zS�Bm������<��?�(�=�T��Ԫ�6����%8HU��A[<N��:�1u�)�i�5�o��[���:n;��h������e����|��(*	��9H\�%��W6't��f{+�;�&�jp�C�ůTt��Bv����#Z�`�V�-���"�g�B����Ԙ�H���rh��X:,�ԩ��l�28��1���8���:=�'4i����[�"A��W,�T1U�'.�i���t�%b�]���^��+cϓӗ$����]Q��R�7+ƙ/��`��^�qBd�����eK�`|]��>f:p�	ȗ/�q8EX�3�mu��y��$��&=�vO5�	��!D9>� ǝ��~���*���ֲ�Q��y`�t %��% 4���u�� ]f�>'��K\JS����",����ܪ�,�Uc�ͼ�N�B�o�<R�*>�/�_�n�8����^*�=RfZ�ٲ�37/'Dv�W\q,0�8zrjc�	eh�43'����rM��)�ߢ���G&4���.����5�>GQ02�N��Ɏ2�R�s�z�C�+���?����\?��Wʹ���"�w�U2�jA��EQ	��|���$Pn|1���ސ"����9�e,l�P=�{�_I!8Y�r�展6BL}��G�W��r<�߲)1Y��	� i���*���a�NU䯐�LY���h��>@�����WC&��ذ�[�s�I�����_�)>�s3�C{j��x�p�]1��J;E���6��<��}�i�����{`;���í=�̇�HK��T�ҷ�z���@�ز�����ciY�I=j7�{�1E�Q�҂�����]G���l�����I��s2u�'!�qI�:2�B�s�u��Q��3�RʻO:����AD��Ǯ�E=/W`7��
JT�M#�K�3~Iv0������V�bj	�͒z�CP��ތ�*�p����g�]r�g8�UY��'_7h}���]p�g�n�ǔs�E�X��V�㕷�X���̦�,�����i@Q/��1n&��[�j���?>b����&1� d]��*>J�����΅%�5x�T�Ov�6w���_�8���L�re&Ӽ슺��53��;��[�ɸ�2��-�"���?�*6�Ա�����1���tQ�Z-v.'�!n������L����1�68�V���T�Εc��%�؜�kڴ=,X���(�-�\#�N�W:�ҝ�p����n&��iy��T� 8�N��Y�y��޽��6���\8)}Ss��T%�)����4����A���%}2G������쀰E�F��9iz��J��BUko��#"�ĉ��\�r�\�s��>�
�	c��	�S��6��ܝ�08�'�Y��p#=����}/`�����sN{��k � ��Nv���L^䎅���_?��zi�;C�n3:�d쁹�S�����XL��g�	����������;u����ͣUZJ�����:�{�S��q4��nG�>��P�/�B�p��W�o�z,p�[���<1)��-zGk��H��_�Q�n=�C�^&Q��a�� �n@aP��1���m�~���������|U��p��Q/1. U��r����Ø�6=�x�x�d�KX�����(8������K�,Ĕ[�!�Xt���G$l 8�E��y��FX)���HG6k�U�o�燡�h�xe4&ce3�}����*����6��-�B�1� DTNOa�,��_�t��cz��/��ޤ��
ȗ�B:�e�-���q���_Q@��UϽ�j��MA�Yٲ�d��<��v���6���1s����s�SQ}��m=�\�X�6�D�|}�ᝒ.�A{p㇏[f=�q�RK 9)"�ƮY
���!��9œ,r�t�}�{Q�r�wP�<l�����u�A�-�����F-x_�r�1�P��0�l���Y���ݛb�ʒ�����'���U���hܬAZ�7�|���Z�u;ZF�]"�,��ɡJ���&u���7ST��?ǌ��Y�u�6�e]���������cf��}x+��s��?���	I^0&�~�� S�G����q��vt���7��.:sIR,�4i�Hbn��GY�m�H�yV��(ܱa��8%��58��͑��{:k`���n$R��w4��Nzr\�>��9��Ѹ3��K���S�u=t$��G$����W�Bd���X��7��޲�h�2��@��r�����ŝ9/���-����s*������>�XJ2�����h�N�&Z�������Q-	�������13�Z�8S��(���8��j��ČuZ�Q���BF����y��G���f7a����N�|��ؓ2��O�I�	�+^7�V�{�V �����v2�<5N����ND�Y(�K���C!ഇ��Ũ+�҈�-���b5�������&��0��3�S8�1��܎��!a��g�'��=P�k�6�4P&�D���\4}T�V�!��pV� /�`�\�%��8��et���J��W��@�����%������u���i�*u�3,s�Pո�@e��Br������C�L4�|m���gEp������e�ա��ѽ�,P�_x��:�mF��2���V3�D��T��.�6	��zXK�.Z��]�ĸ��2�����ޘg�o0d�:������eN�H�#N�Ir��ӘF�T�D��|H�Bַ�Vg�1���҆S0��pC2��<sCF�� ͧE?�Byp�v5��-f�mP.�*!;1`NF�0I�(�a�*�|+Eg�=�c���6���:{��j��y�����O�_v̂v�ES�;B1�%ہ�}�g �P��G��%Y=����:�V��ʻ`�͌�K�.rY�D�}Ք�>f;��{y���H,������4�KF�ӻW����[���m��+�9q����)X1�
�r���R�T���dg٢�7��?��mb!ה#�Hd����guX�Rq����ھv�6�#ö��/��S�uw�T��ח��b?��W1D��hb%?�D���,����G�~'"2,��X�N����+i�fefCnӃ�{[=�9�D��//��]��S�h�D�]�"I���Eb^y�ٔ��7/K

/�Z2��'��1�3xvfP�#F��3��o�2&hr�G՗Ӥ��|%�˷��!db�ŋ�Au��SoBX�������D���%� ���{J��-f��{�5��{7!�Wt߯Fp���������h�~rz��Љd�Q��}'��4?A7~ ���"��'p��5��Xەp�I��6q�X]퟽�0NոH��k�pd&�2���ۚ9t/��8��k�r7G��]��jv��	8DK�x�=�sJP��֕�VJ��&=	���E���~+0Ҡ!�U�*@9���&�T:o�3�����"�K�G�*u-,yBW�Jlxo:�: DUjZ�GK�B�O���<	A�����Kݤ�����60�'�����]G�k�T@��@qY<�]����w��w-�7�|�M1f���2�k�Lű�Ď�6�������~�0;BU��)��;��G*�Gc����'��D�d�sO�y&���?��*U�[���wp�	 [!)��#T�:�6jJ��"�oe�����n$��#v�4v8��c�=22��[g�s���/�r=��[6�K$!j9^����C�w1���IQ�D�RK7R������З��<X"��Wh�x�h�I�`+�9W����mI��P�u��	�;���D��˞
A�J�@��ø�k�����v�^��6�@<�ϯÿ�M�%Vֳ"lˀC*��pY/�Ћ.8��QwpM�%U�?ц��t"_&�Ѻ�J.�}��d �t�)���N�fNӜ��ʎ�9DP4+�:৖�\_;�%�EAS�� ������N�YR����_*���j�`�l���4�V�a̱��-�^��'D��"{���;O'�u�0�x-i���`�HL�N��lO��M�m_7�}z�w�@�7	 -#�����9f�#��k�`��9dq}f���7�_ Iy�!�^w���md^��35qMuЧ��	~�YP�̒�f>����Z� �xk��i@1��|��X���]�ǔ�i�9�h�S�RZ+dz��4f��2�8�?6����wq�c���60�c����[gL�r/�.v�1�+)R�db'��	7��֥�pW}p��&��������E'�+e®�t'��3"\�4ӸZB�|��"J,�ǭ��X�$ݓ�:���&%�I��]:��h�`��k�3���PPkN,�Z�îᾞ�5cRԲ���#^�y�����׉! 
��%1zҝ7���S�]D~����:���$��O2	��ҥr��*,�x�1���V���{���=��E�7��M�h�R�>�W�ajQڀ:͗�9���Q���?c�ͧ�,`З=�sD���м�+�����"E�
����D ���0�܃䌗�Y�w�׈J��r%�hb�]��4c�c��u��s�[�JD�ɛ��4O
n�?��~q��^���j�/z�r�;w#=�n�~t �<�fٽgct�e�>�\UT��1�f(�RH�(��Ƶ8��"k�W�D=�*�W��֢�T��a�+@3�hels��VX�b�MFk�� ��#�������
�VeUQ���!l�%u����'s�7_���2���9Fм$v@�@�K�0P{����-�"�@fF�a�N8�y@�.�i��չ�Sb�ʓ�K @�kْk���F�I !n����6���JHk]Q��~�f5��&J'\A��r�:w�y����tL/��̪��Tt��<���:S��:��e6��L�D�� (ɪо�@?�$M�&�<���g�16�b/���ηO�-��:+��%���2|�����JE���'�3 ��2��o����3�(�a�v~�z�1ļ��(#�O<����.Oґ1C����p�C��(G@t������ C���2Z���2jlX��d�	�-���g���x�eK��\�ݷc/�&v�ѡd�Z��%�*�ֹ$5��F/�"o��Ժ�8����P�_
���r�*0�N=��7�\m�mI�gK@��.��~��ji�� �hn�'3ʻςcчѰv���wjͬ�n�А'�V�xu��W�F_�����E۩Aoo�	BTk5}Z�����	=�ʒ�	�sx�5e������9L���~z/w7�k#T-���8B��R[��>�ۜ$��^��.Tu���&�}8�7�E<�׻���Ɏm\oQ�5���N��<g.6W%n��\�$=���㕫�PЇ�P���Js!�7�;���V��]���%���#�Ġ�*~S��!���M��Ns��M�f<ܐ�{)T�"��%�� �#�9��*LT��fV��<NҸI�����WhԖ"b[�1D�˻cS̚:��|U�KX�u9����GP/m1M�0.�vUFG�Yu�\�c(J"�׫"���s1bq]��CKa�������%���������v�2��?l9_�['I���P��K�N'�&�ʑ9���n��\!�<L�!u��%p�^/y��j�^å�o$�"�-�-�y(]�\ԃp?�3Q�	�����r,��2"2����Ջ:��]�_QpaT�PXq*�*S�tv���v��u��������6�c�&wd��9lN�5�A]��� ����_���ڕ��mO�xЛ�������)5w��h�Rw����K�R�IGF3�!�B�du� �Hr�e�NN1=36�4l��1��(�{���c� M�&G��ߌMG����t���_q�;_5��N��7�&d��3t#�4�C�}46��0Vz�;KiO?����M��ƫ^���c�����J��v.Z��3�t�����e��@�"�f������I�ޣB��6��"+��r���Q�L�@���s��'��.��昣C�+��c�΀�����|���@0H����� ����}�!+���vó1���d
��]�]�y��響U�� 1ã,JE<�V�´f�jټ��j���xېpM�W6P�I�Si7 �T���
�j����{���L�ӈ���5�&� �07�TA�v����WF��8�i�p���׭��|�t��ɿ^Z5p�Ώ����V�ʆ���NP��L"Yg�9��oP{�J���=F{$Nu[���1��~h��4E4w�m���6ܮ9� �H���?t��p�a��Ƽit�hf|np��%u����4�W{�A�8�b�ֲ�����RȽ�fmq>I�j�!t�&���{59 }-�Ƽ��b��?��]�����3�+�_��al���Ն�7�a���2HT�NrI�%�.Är�G+Se˩��f,�t�f2�|�]R��;�Ύ�9>n�̡tNl�оi0�h B�3Y�n���61��\<��3NȧIz���t���H=hi}�5�h���S>��֬�<B$GiO�\t��o;���M4GT%~����"�;W����cc:2�KXZX�r9�\q�]m/%�"H?N�e9�wU�L���"���|��/�.l�qF�᠊6��q�<�N}�> v�S��D�r�f�l�:�P�����҄�]���%�-�
I���Ӫ��/[�c��U��
��L�Iۂkqi"���sz����A�I�r)�>�G�rn�Fvv}�wi��JHa#����d2�pk�G{�Y���3)L9tн|�>	zEˡh�Ȅ!�&��i�~���&�ъ,��-/{�B�\[@��6��ۻu��^���RDȁAB�f��s�S��H&/��	�\6U��Q$y\p�߽�7Sl�}��R�`a�davL��}l�Asq]z�&��]�*�ϣO;�Z�_���=D"�e3�g2۟c�	
3��T�;I��,���:)q��aZ7eQ��b�lmN}�����,�;�϶^{���s% i�����8�Nϰ_�W}p��0�f��o�%�I�n�x��^����w�I��"TM�3�_��|��c�SҊ��V�m��$���-�`��F�z�V��z��T�#ʡ.�L�g�[Ljj��ʊ�C��
�����0���>I1�息�����F{��6r�s8��`'���#����yhQ�[�Q���	X����5�2`�w�
����I�R�۷g�>��(�%�?�Hfd�߷��7�e"|��~p}�R3�(��1�x�۫�ɇ���S$���j�<Eb)l�>-�[��6 �*q��;���i���SR����P�V7�=2ú���A���P??}+����Ʈ�X���0v�ʁ <�|#vT�;�!8��L�ޫ��za[H���<����ks���ܱ�?G�E�="6�}�+w�鱭T׌��*���ȭu��,�j")P��{�B�Ӳi�D9�뇎$U��4�:�iJz�/#YLU�ƞ+�f��r�-\�y�Hr��g8���9'��o}M5"Tw��c%,_Аp.�@�j"��3�1�SK(m�3א����\D�*�#�g6�G���Ay`i���pH ���	^��|���sp�W��4N5y�δy��$���ؐNm -�-;WIx��K�>�@�!�)�����$ �<�Y���?dw�K�.g1���ɍ�P��
�v�?�$�6)f�F%�Ua	c=6����hNo����+A��r*T�+]�u�H��0�W�뚗-q�W�|��J��c��˻Fk��ާ�ynj�A%���4)���>�Y��4�l'��Jc�!iR�=GK�@�6b"4�(�`0h��ar�ۣ�(S{.��_��)ռ�?-BC���]�@��|me�GO/#�kuG�ڊ�u������*��]�s�c�jy���ζ�!Aۖ'�Gv=~��_�_봺�h�<�c�:02�A^b�!��|��R}�`P�_Y���{��,�b9,{�&�_�nls�6�X��?����ۂ�@��2�TN�B�/��`�8�t0��e�8��ո�C`g!H��܅�TJ��c*N5�{���S��lC�ţu\�y:�3�t��'��	��S�k��J	²B��G3���� ��8eq94�i\6-ݾ],��.�4}| �,�I���x���􌎜����c���u1b�x� qHӱ�o&%�Q�Xe۳}�	���Mae���S�`_?�~��
�������������M�ط��U}�#�����@���&Z3k�`��3�#�x}V��O���0����&�8���1���Yl9��R7�}��aE�G�k����b��rw�k���ԓm5������T�w�G�U[$��&�+ӡT����;>[O@{�f;�����_*����?͹��Z�]���k��)Sʔ��'�=e[�6eڬӋ��s �/YD~^�����Y��+д�C%��7GW�ڱYT������1>Y;,M4b��fAT�xJ�޲s"���?'"��1pƀ�d�[%	��~�G�7q�L�2��e�ܛ����:�gQ�ܕ��;��A6_���gYAl�ì���h��v;V��n%H�h4�����$c�fV�����[�~�������YF���HU�+�wCN$�����3ѝ��z��ax��}Q����:�H��aGi���!q�����߲�������{���7K�]|[������'�<%f�%�v��V�\�Gc���A��K�Ne�%ICTz��������/� ��%��+��-���Ѱ�csi&NȢ���VpD��s,OWu�懌^�������-�,u�mdy�H�[�7��} x̢yVf?��n��geno%]&N�e8'g(�����}m�3p�b�s"baG2�u~��8�sn/#���h,��į����@����Б�k|4Z����j�gu|S;RK�l��+k`<͔���7��M�i�~~��Ko��Ui��zl�A������2DqҐ�1��c��?��'�}��p��$P�偅�d��1��ԏ���ӦL�1����I��3�W����@�33=�i�2]Y`@���0�fS��IXw�F�E��N�(�jo�Xk�R_$�$r�tF�[�7�� ����Q��㐽�uo�Zl<~S��$��}H�ר^?�$�u�]>CD"����Xm��5c`��
<�)��g���a����%ƚ=(��r�֢[e.ƆSnQM�*�����p�JY}��{���&��1��rD���Bިۊ>�1�
J��pU"�X4a���{��a������q�����]�GD��%���D_��'ͅ;�\V��*H#:�F�$o%V��Hy��8Y��
Y6�H�s�<z:��I��L�2�z� ��M4��޶�F�c��HY�G ����]Q����@0�B�{O#�}�a�Rh���=#}����%~�@�?Df"��t
��*b���N���X3{��B<ܜ��Yfϻn�b��0���*��jE���=E�T3Rc5��Ȼ��bS��#�����dpFq�X�S\��C6[�CJ�.�Z'o�݁�PK��fS ��Ƿ��Y����=~� �����au��H�S�A�G�d�p�W_m����Oư&/���D���~��%1G��E��.�����+0�+9B;ő��!��Z��\�.F��c�ݞ���#��h�˼o}K���8l�P6v;��j:�:�ի�����x~m.�����yl�NIv�?�
N w��
�q�JG��S5qN)���Y�m���Ac�	�L���p��D����E����F���S�讲�/yú`g�r���5���)�ӘS�y�6�J�ӼS�tg���N!@7ԕ�Erl��J>���^f�0�h�Y��
�OSYk���W��S�n��Ds��z�`><���Xl�����RQ\2	��}���+���|+�Ua��`\4�Ff�f�8A��M�I:EOMH�`{��6 	�&�2��X�YM25�����!"�73�s]�E����2��F�y=���x�}c�ݞ�d$��>g�)�6> �$��k�
 �=RE/Lf����  t��?���t�� s��6e_hҧ\`F_NMaau��NeɇR)P�S��$e�<��5t �)�(���+^si�9b�<������4N�%i�#S�1��� bY]�N�7E6>��~��s
1�M<��[���H�Ά�Ă�.׀�/y8�rr��c���{W�`47�v�r5ڧ��F�!����L����ȃ$'^!/<i�T��@C��/�Q�5#��>�^�����Ӽ��d	]�ӏ�LϺ>��^4aL�N�z�|W���tOGh���O�li@�tB�<��\�
?��c~�tf[`w���ʯMpk�w�(���ls�Qe�{�d��ū���p*�ФyRg:f��w�1 YJ��O.��y"�u��)��[?1�٨��}8҅�Ŕ$u��Ono�ċ,�Hð�a� �z��f"5Z�*��4N�y�M@����T܎��~��s��q*���V2�/ ��T�c���5^�x��
�G{l���K��DL�k�n1� �@�,��`���M򅕖2��b%�x�z�y@�KԐ[Q�K�߁4�FT������**��Þ$�����f�,��$�A��&����;<�hq�L��d���K�;�f�GP�6�Ů�"��:�������w����ݤ�8^���ό?&��������z��)��� 6v��]*n���ģ�S���_��B�a�y+@]��a�	�����t�N襽YD���]�%��%��2��:�6jG�6��Gqv���3�zkQ����z����Z\��ܘ��n�*[�-��g��q�a�O�F���м}��W��5�n�>�H��0kRݞ[�G�̍~X^6�m6�9!�v�����o���>��/��������w����M<�������[�X��G W���K�����_ >W���:����핛�9�Bܾ}8)xtr��c%*���� h���ށJ�_�7�`��z'Że�����8��Z ����ٴs���_Zdc/��6������-���n�����N��W�,��&�#6�?��o<���}��c���b�5��ϟ`ɗ.)�'��	����L��<�B��ʦJ�n� m���)�+��w�OU|�1	��ڃ�c50]*⢊�AR�}���[��f<�R���g�	����BMu#��K�J��#��&Y�����C$2�攨��D�;��v�2%1�������n2� �`���=�ʏ��P��CyM�\�^�s�3�/0�[&Q��<���2(�>=6��j*E�
�J��h.m	��eH�̖
u�O�Y�I����-BB��|�s_�p�Z8��W�Tc?��^j����s{��9&�r���vq��	b�J��5����͑J1K�����W�G���Ϝ�jz�Q��Q _�G��M�>�X�4��.��p��֎���e'#s�}k�u"H��`U���ĶJ,�����W�kl����LŢ�f�m��2�6���f���{XK�J��A��`���Ua ���7���\���4,����|IbV��� O7�i�Ow��nhJ���j�Hy��@��r�Pcl_9?$��oǺ�>׏��P�aG����&����4�ٺ2��h��l�������p�:����U�1a�� k�,��"I�f:]���v��K���+|AU2{��&n����|z�u*/�޵�~�P8r#.���-ȔP9?�7�;�ӞH+O�b��㱡ė`4�A���]x@&~�s5�����'�_@
a|�@�;�j�x�WS�q��iG�c{��\��@/*JKQ��*\�ǎփ�2��AG
�Ӝ؂���Q:%��2���`(	p�.\5��/gV�C�Ч������Y��)�X��';Tv`�{�i����#���jr
� 1(���-}7����z�ֆB|�ĺ[8?�z�4�X_4���I&�ӿ���b�)�hӧ��l�\]\UIrs�WwrQ"G_b1����PY7-Q�*l�1v��=�Ǳ�i'����Q�� �!�a�|�s7��<��4�^��P�!h4���3�R�׺6�\�ꄒ��::Å�Ś,��н���NM�'z����1����5��s�ӢMѮ��9gĸ������V��n��f���4������?D܋^'�$��sb�ц�κ��D��쎂뾪}�Ҿ!�ͽֵ��-���1x"m�_�4x���j�	.g��b�vs�q̞�Z�u�x��x�d��:��ߧf'��ĺ3N�������q�=�*J� ��bo���!�ڲ��ׇg�кr���dX��)���Yu�r51�3ߜ��1z�x*wY� �l`��oPI6�3Q��|q��o�OL�ӑ�折u)'�f\2E��P!��`��]Q{��֊�]���ہ�����ἀ�^��K�/�Զ#t5�I�9��k\h�����0;�xh!t'�9v���?oH-"����-G\`�,j�F
�5V�������W�x���|	�0�2����N|~&��x�P�F^�u��c
��M5�ZI��ۛ�@�G��� �����t�*{��}ܼvA��D�3))>W�c{p}�� t�\����t{���^B	�%Y�e|12%N�+���IB�=��\
>-��	&�ڃ�^�p�>�*������`7;�S�e=���j�xTQ�.*���<���e�(�@Ia�:�٩���"�4XMD+(�$_��;w(YW��`�M�V� �?��z��)J/����-�5��z���!	�qv��	b��b&�����N��I_��U�D\w����rs��X�����������8u�96i,[�\�@G֖"E���yP�d	h�t���=��:��g���jo���a�s5�(���]�A5�邔��I��(����r�|-��i�ה~�/$�Rߢ IYRs�u��n�Vs�u�~)d!J������-!��e�.߈�M2I��W<��!/���lSeH%�w�?�x���͘4D�a�M��b֢Ȟ����f�aR.3����R�B��}��=�&�j���+s_v`J=K_䄙��h�Mpŷ��O��y��-䦢������w}I:�Ϩ�r멂+��*�ĽǜWڨ^�cŞu������2<�קҾqR1Q����f��ƶ�(-��lh���ދ�p㋃��;-=�o�L`jS�}՟�&���cP?����3�#�K��_���_���8��1w?G�\�����)ΣDB����O�-��~� +i�F�S3���\}@����VT�Noa�TGO�`2���F[�T*�
�ld*�2��sT�cg�^ݜ�׳s�|�2�̖��2���MV4�4�P�;�q�b�ȿd/:\ ��?ЏλF��C��:.ɍ��\0�z�BV���@RG�U��Fۙ#�Ƿfu{�m���1ic����gzP'jF���%`�K"L��c�6�?�{@�j�q�8��88x��:���(Q)�����T<p�՟����D��^Wg����h���)��РZ%�^!��@:�1%���y���5�8?v�C9+�Q�2
:��7n�Mn4�|�nU OU8���֫�V�&a�.��Ɛ�͊Ex	)@ #��4RՖg�L@�}�wm���PxB�Dg�֮�f�ݻ��-�
mt��V��n{�*a#�k�HGq=t���3�F
7> 0�;@q 'e�#��g{5_x�UTI`�-BxI�����9���E# cJ��N��/�{����}�Z"�l�M��H.�/�
�E w(^:�;��u[����{������<]{�ʺiʫBIz~n�ԁ6ɸ�	�33|�8R�D�m��3���~1�a�l����7�>S�Ј��cC6�iӴ�&����Iq�뇀�G#D��=�Œ�E2$gl���B$rX�g�Tt�R�[������%	���|c
���-�
a�ᢰ`��s�	
1=G���=���Jy-55T�ӽ;��$���ez�4�`��[,�q��T�����JIu�q�ҳخ79r�i�<ߊ�����
_�(�+`���n��ME�Ua�٢ϫ�1���$�.݅�~{�B^*9�����ɛ�d��Z	��_�	$����ݺ���;���Яz�	}F�㯪��C�i�mXG���k�g<�݌� ޅ�r�;�[_�n�:�u����I��Qd���G1����k���H�`Z]T~O
ݙ���^(V�H�TK��OS�@�F�#��m�ñ�u�y$��Vc����9��m[����ͣ�9�e��Ib��?ä�o#!���C�Ƴ/��)�vm�\^2d�9�~���eef��-"� ��/]��T�aT���E��,�n&4�:c��㡟��%Y[y��;\�Cc�;�+P3:��9q_�A�#��8Ȣ'L��ڍ	CS�-�x�DPpG���©)-�]���JQn�#G��S��|��t���
�`V�V\��4���{��÷�FA(�R� �%�]L�Xh~�1��p�>.���P�r�E���v��k(�XJ�i]JZ��!fۍ����E��0ק�����������1iM�TS ��;�(C�P�k�!�߁/���
���T�_�ݽ�
�C!�X�z�$�]Fv(�ݶٰ+�F�<�7�8߇L����I�JYd��zhq�'���B0O��������'�t�V黬fV�tj��Wi�����p��{^;;�iK<>�y��M��� O��
l��;���7���N��5�����n�ޓ�H��@Z��e%�c�.]F�pО3�!�M+J���5�*��g��^+�"����.Ԧ�[��CU������Ƙ�F��gEw;��G��h5��U&O�4ojy�Ҳ	�x���Ŗ.3��͚�ݛzb��1\��ْ�舾�����o��ʀi �]�c�@z6IH]���і���<�'!��S`_��`�!��1���Q]"R���[ ��R�5O�6����Q��	�E�3G�n��e ���n�����!��H����4��D]�<���d�G�J )���3$j�ʇ$$0�Ц�l��@�,~0�P56[R�����yrI$I�h�ƊD�^Zy#���z�/;/���Zu)}�@��z�d�w7nӷ�P���b{��']�sH�P��� 8>�rU�mϠR��
V��Rh�.PE��b���z�P� ����|>h�*���bӯݿ�D��� ǝ/�^���BU���B|�Q�g	 v�,�;&�C�(��q�
�6]o�Q���̖z��V��V�Z�bh���^��c�;;�.�R&~!�������&��E�Q�G��D�P��B�A�����[�|%(l���Px�x�r���%>(&'L��b*��>c}�J��c����cr~�ؑ3�h�y�ZW
��|�L�@ ��Q
�!`�5��"oe~��\��c)��E�,��������l�A~VQ
��٣A�x���A����n� �AD�0yD� �:3��'�a��D�Z��J����w�l�:�+OgL�S�Xo��(��Z�v��=��\�:} �G�,f�yh��8�a�#��%�/x����}E�֙�ê�_����������7<�0I!�ә�lL	�+[J^�7,�i8�!�7"������F�)�� ��3����+���"�ܳ<�L$.-��6H�N�Cv�/"�l�V6RA�:#�FQ�I'�̣��I�k>����<�x,˾�O��9��J����~�-�w�����&&s�e�����7��Ԏ��Xk�y8�3 ZJB
�����_��~n���8�6��I����a8E �?K�Cm?�^�r+���c%"{RȀ���%�ړR.u6�摌7�>�����$~�go�ng����1����U��p���s�bL��W��sp�ᮈ��g���&�#��OmL�.�����q:D I��jCvpk�/@�K�0���3���צ��ۜr4�m�a䷑��1��S�ۄ��L%�?�Z�����w��n�]F1F�ٜ��8��x��KN����ۮ��{k]bDd]HYW�-�b�sM��P��m��u�T?{{ng�;�A�i>(�?^��	��6e�1WٱN��Kg*��j+���D��["���dҿ�x�v�����]N��lv�g-U5*�<Zu-b<e�.��h�ޕ����Tݨ��ꠞB�A�{_#GBQ�k_<��R�gkC�L\�Դ;����(:��[J��Z>j����xu;�k+� Q�Y��Y�����5<G��#����L�Ř}�����,��-� 3V}�R�J�
������qDGs���a��αiYV��@*�������Ѹچ]i�U�%��	a����jʁ�M�-c_�\�Hf�ә��P�T��$�45/�v������i�΀[�M]����#�T��k�FމЭx���?<y��KvH�Q^�/Q2U�a-�fN��YEg.�����w�#oz��Q���R���t��H��C�'�};�yh��]�D�S���{֜Y/�9YR-CJ�2��U�q����Z̷
e|_�y��~�U����f]0���� S�l*��h(�b�T�snm:��}�*�d��v9�y]�R�s(�k��3v?A
3͜YCG�L�UŐiP8v��_�0���B��ȏ�(X| �y��Wy�k6�nܸ�7�SH.�f�5<��[��ݤ�.�
������쀌�g�O�풇�ej2��pAh��ʚ�y��^'�+��P*�R�#^ @c�2u�r3@q9�2РHI;�jC�3�DHm\[_c<�&��Ă)�<;aM�L�4� ^�[Y�����RpE����4�ʝ�����}�d~��IRQ�� (��CZq�lƓ(��Ud\�b%��6]5T���Tt(����10iz{�aN��}t�d�j*�=�I���>������|�����[�A��`���k��Ѓ���0�)�v��y1:M.n�=����
*sH�M���7�N3ȧ�[ rR��b�29�fZ�ϲ[p;,Ky�הf��B���l��c<��%����T��&ls��$���mZ\oN��~�[&��&r�z�p�ag��+s>�4�z��ْ����Hxc���
\�cID�
c ��<�*��͐Rn���е	>_B.4�6N�3��=)�{���t*b��DJ���u��ɱ.:0�ҭ<oj��2Yk�L��f�>��g��� 2v��3��v4��hN�2�9qAŠ�����tj�>���b=���a�i�q��h/N��k���d3��v4���E��`����o������qh��?�P��6���4;�q&���6ֹ-��]ąDPN-q�r"�}�[�P ��g�:���N�
͊�"�W9����Z��%��qq��⚅%������)��@�4�	ϢΉ�Zr�=�%`m͊(g��{�� pS�c�JQ,����`����0�����;?��UR��20�+؋�桥ke���1芀@:>��Nw���ؑs��c�f�'��k$�;E�#}����:!f�}����3
w_�jn��!���C1@����2%	�,�q(2�h��!������$X��$n��^I1C�0DE�N;���ƠK�����+��uPW'��{Gm$Sj]NQF�؅�R7^����(1~~�E���9�f�KO�k0zY�v4��?R�9�OU�Y�5[㘦}g���Xlp���Q�\֝Ѵ��:�fIM�p�C۷�b�Zo�Rh��#�~U%`�T�y�kFO� H��h���+�|��N�s�A���y6�Ɛ�CM�bf�k�Q�H�����{t�.�>f�-F��a�Xovm�ounP>)�#]#1��ɟ���r��Q'�!N�Z��	��9�N��?`�-kp�˿7µ���M�F��~v��$K)!��ee��e�	p�p4�(�h�7�D�us�J�U(����.����^dͿ�����K@����\����r��c��K}������d�3)ߐ5#�+!@��E�de�&�W���G��������"�P/ܝ���P>J0.��D1���XG����$�`Vd�\&
D�� �&w?���/Jh�ZS(�SB���LG�B�(�^�	"^�T�(��A��N�m����1�V�G'Ձ������2N�t�G]��F�7":yЦ��#�Y7;�RH?o>�|xP8���@g�;�M4��vO��(�߻�m�h��- ���-o����ghWK� a�[�7ep^Ձ�q�t��ڱZ�A��h��S��7�V�uE�b�k��e=��BYK(�-��7ۦ2i��aG�l��a#+�Jh���)n	�4�ʂ��a�{�wt��>	�m��wY)�Ž'E �U��o�$'��$t0���c��@°��/��t�����c��i�����l@�qǳ����Y{5 K�  1i2i)���/���	ڔ�䟴
��;���)^���柦���,U��y�zd1"�MT��;*�����������)1�9���%$1���E���>S>���D�KJx�:v� �ܡl�����'*i��!V���.��-)�U��2�F�/`�m�xÙ�v�oWJF٥���W:*��1�hDR �~�R�5]��>gd/X\��H��E�v�̲y�WC��F����#��+R���B Z�%H�yv"6�i��A�:��Fg溪0&�F�[�1L���	��F����1'�Ć��n/T9�pᰑ�=���U����Á�N}��s�%;pNy��]�s�ǖ�e���/1�C�%�Ky�c���7�K1�p�q,<�#��3״�8���"�):� ���ym�s�0��ʇ�T�~�SR���w�Ve��k���ǒ����$l��I�@C>�p���n��頟�&����i�U�Wf�i0>�۲?_��v�J`?K�������O�u�{C�նۮ�|���0@UG	��W��d��`]�)���3'�XK{'��x,�.n�t�CX*��T����ȫ�4M=�p6��b��:=���5^D�;
Z�ߚ��.;`�jC Vjf���2��?O��ٞ&>���!�K�B��������9|�W{L��� �갂�к|͑�f��-��lY��P=Xyx��0��.�������O6X�Z�ϙ"(�>A�X�mکHG���k�}�\��0�T�$Šo�M:�ZU��
�L(/`�o�Ķ0�>�^�w;�q��lN]�L�*p��}/��:L(�Hr^_} �&솔�'1�(,��Ȅ�o^�;�X	UY^��
'�*����L�&�Ro��n%�ޔ�H���t���\�a?`�$�3�,B�_��G��&{IՓbΜ��pHe�h[6qp@)?�N,����pB�Y3b-�+���z����v��K��̇��r�[>%�y2�*����%1
��1��~���S�Z�vV;ݙٞg��t)B\ɩ�"gtsh����mqY���'���#Eη�>J?���P���cI��.4�>�=���W�37gkLkA߰��
�>�{���f���D�4
,��)���T �q���0�zه����zG~}��Y ���p����V��pH�����!�9�^"��$���4�k2�`D\�H��~�:��!*�`+�p����t��ǂ-QP�W[�Z/E���e\����a�C�k"/�'\��ϪH�(�|&��̭�(����V��O���F,�0�J+�<#�Z��-\ߒ.��y^�
Nr������=�LgY˝�>[^p��0J)��*(�F���W���K�e���EČ ��1 OM�%J��T��׾��z�7)�m#���]W=�=�;�[��!
����΁r!;7s�qXuc�$��@D}���f�cBA?o���[����:qtU���l�=���?řek449�TqKS����I)�1��9av���]ǟ��@��%k^��l�IOc�D��]��Y������@�U&]����d��_�@�gzV78]rf&9��Z<T:�����=Rg�>r�Xt�|�����Q�<��Q��-r���k����;O�=��^nm�chY*T��?W	9��*0`��1����0�U�/<��8͞�5f{rH��4�C��#�i�)x�!L,�͍��S�O�7b��s��P��w��៴J=���«�:�k���8�:�� �K5��F�\����]��D���0�ڀ઼�˘E�g��V,IV'���ϓޚ�1<.��#2�
�o�<����ܥZ��mp����]����f��<��ޟV�1p �s\�6a࿇�e4��ZJj6���1��r��b��������7ڬ�b@ߚ���q��Q�8+��T�t6��M�������0fd�N'7G�����s��v��'%ז!gr�C�	St�剰����a��Ǭ3YI���q�.���҇#go�y���U��Yo46�\�T�2XyG�m4���Sr��I���S���#������&c%�t�<f�+F;���E�M��}�_�~:=o9as��A��!g�@#?��q�~d��=h����&^=X�ڜo`C��륬��vƸ bi��Kp����^��  adoG"p�z����D��&��0���ǎ��;���g�AnBtb���q� o��ΖNE��C�=)����ErY;;&e%�g�˯6B���oǤ/��T�˶QA��"�ɺ���t����	/��[��F�ɥ��Z0�k��y��CQ:��%��ع� O��q�n�������nDZxjm�����~=��2E��A� �H�?���Pi�mU���}y�6b�uz�{v����t^ڥçr�PAp���L�c��F�F�Y�ΐ�0L�2����x�ͩ�iZx��4�}���6�(Su�)�$���򐳿�V8	�����P�s�QgU]�Mۯ��ןQJ�6,HR�G���2Wu�/�*X�9�txLp8oA��~kp������4_]3�g^H-�Z
OMS ,���-/\1{�L�?:J�����z�4��Q��%W�DM2�G;��s�n92>Y�p��?���,�y�]������M��z~^_~M�E�B��:G~hIGq�F\-m)�D������UH@ӎ<
����h�XX��u�w��~Ͼ�Y/ѳ�]�"�v�8�hW�j1��	b�b��_ ��^-��ZЫk���^p`S��)��Q��K0��ɮ�sO4�����y����-N�n�+�X��\M&b�X�f�ǌL,p�1�Є�8�g��:��l�EK��5�/�.x�s���a�Q#U�K#bg`t���S�I�n8(�F�<@��w髙�h���/Q����u,<�@s���e���'�d������rѥ���oՑn��C���jL�,�A���Q%�� �9�V�8��{�8OCCIe=���~9�߿iaXs�$d+��^��q
�8 0+�|o�J��Q���+{��(cf��]�Ȱ�!N��4�BЋ��HVW\,7������9�0��~�\����@{����#G�N'~7_"~e}����~����>脙Cyv%���(FAC��"aŨ�߲l��[��%�W��P7^�%�,��.��J����P/wƇ"_/�(.L��[��4k�uf���L�W<�֛�ӕ�Sk�J8I!}c����+�b� F
���h�]�������7����n-i96*ڿ<�+U��+D� c�o���a�U��n���ټ�U>sjyǾ(+��L;��Zt��$,��A$HE���i����>�W�abt�X��%yw���z��A�ʪ�18@��{:S�)�+]#���q|u�� g�L?��E�W�>
��I+�p�!upl�u���I*� �z=�-7:E�E��G�꼫`�IY�ˊ��p�����������〳qe�!�z�i�XS��f�	�=pvh��ĝ���\��_�S%sL�U���C��a��-E��D�X����4�'���D�G�%��7j+\&'F�&�!��ieO��l��xJ㈽z��_.����ˎ��.�˅k�>9F���rۛ�ߪ�8F�'�Oο���O)*"��;��}����1����9޷�Gޯ}Ώ��c-N���E+�����~���&,?|���g1v;^N%�<=�x�ъZ��r'��a�P�3�Pr��ܴ
��&�A�l�����_S�m�R�_���[�Qj�����K�7���
�Cs���FXG���� ����/NlU9=�K���a-f���Pe�6z�$�&c|�iC[6�n´(�o����TUh+}����b��:vdk���m��Kd_2D�O��1�]�h|���됵�O~��F� ��T�W8�K=�Q��s'�8D�s�*����gDle�'��j?37��~���{u�"��8�7Wa]��qT!F��T�؏sfm��	�@U�.�����0AQޤz�$a��M�;Q������-;=��=�]7�Zw�0$���'��[�Z�$wl���7I�4-�hSo�h��mQ�fE���xl�r8�v W�)y��;��d8���N?���$�H���h��q��e���x34!SPM�����qĒh��Bg@ ���l���W��xꡘ�-�',Š8��G��s�"�#���t2���-�"��ӄ��Uq�,<5˦��L{�Х��g.[	M^4���4J@�X~g�����WB	R�xb��jԧ��,�.��oŹ�]�?NB��Q�rӉ���Ź�*���#0Qj��-Jc�#v����&��ళ�	u}�pEWSch�U���%��H�%��z�~�� b�n㏜5I�+�ѻW%�Y.m�Z]���6Y+��de��.������)�#�ۏ(^W�:s������i�bĮ/ξ/���t��ү_�~e���:�.���K+Թ�R�Eﲋ�96��(����:;��q���"S��d��}0��
�y�l9~� ]Gz;Ͷu�i�(����JTٌ}�ؼwS�x��2�|�4ji��E���1f�.X�dx�̎�7�7�t �|f�Ľ+9�<]�^%�?�$���f��Q]�g��V_�TZ�)������A�����e[!�I����T�!�T�,���KH1j��0�+H,v�roۜ�(s��Z�q�y��mU25����L	.�a��&�{������QJ����\��B>�$��Ϳl�Dd^u�T�j+���ݼ�%�c�{�����`fn�.-
I�o.T��x�pESs� !��a��&+���4^�b���Ƀ�|���(��+&�R ��YK��<2>���_]�S7��O���d�֔�Έr�7��'�H �#����`S�C�'>�~�<f���Gr�#G��i�y�Aa,���WZ���|������7�<sP����&����ơ>j��̬���_eJ��˥3�{�_��Rx'6��:䲦�w3,��*�s��6��͵>��<���Rwj�]%`?f��=5Dh�1^=ס9Zp ���a�t5K������u.S��0���������7� #�Ps���z�n~m5艠^ۼ/����a��I�\K��U���[�5�,�O�~�A������3Hx:lW4#6>z_�� [��潧����a��g�v��Λ�Y���x%6�(����<�����˫r�N�mS6��}r���NU�ʩGU�s�Ԗ��(e��X��_	<�Ŋ�r�F�����}1 �1[�ժ*=������63��T9UY@ϖ*��b�$Ÿ{����ٺ5���/	�!,\O֞��{����8�D��GȥĆ1�xu��`Ag�gU�R�3�4=���=V�J=�{"�t�������>F��HH?��;~Z5�;跧��U��,�3F��%o�c��_!��o��cU�E$Q�6݇0�pi/p�ϡfb��x�"�.߫ʥ"�@2漸t�v#�b������d��ǟ��8M����f���`��J%�y��	w���~����l���mJ�q���t7��)��*t��=KKfZ��G!%�R�I� $����*�ϼ����
��3n��&�~*8p��@��!4�l�Xg
d�E&��:�L�*C�롱dmB���Hr�T��)��N�E�k�'uW�U�H��C�]�m���3\�L��l��a�-:����FԴ�)IeÒ>P������T2�����O6�(R�����>V��C����O��FI���n��{QH�E&�=�A�`��H���}f�?�w`��o�������c�\Y�|d�)<k��E!%�La�+(	�;[V��s��H�*��N�hp����d�]0-�����X=��U=�,�%�V7�t@G/yr����(5�2&���p�UQ�h��E{9��#����m��z�ty��o9����nY5�(V;�3���ʭ]ȓ��H�boC����>�����^A1��$Z�1k�����I����cvcv�/��sZ��x��� �iDk�)ЅIA��A��ߧ� D��dyƮ��+J�or���b~|�kG��x����X���gG����D�ҟ�{�G��Z>N��~lxl�k5M,d|�t3�	����#��6F��ޟ�wU���i�	���%��ݣ̅�4wlK�R�)Es��u�pO��^�.%�5�v2��KSp�r	�[�]�=g-?�n��J��u�����������Ĉ�u1s`7�>�^��n&�(F37{��[�2���L�U�Fl뇥���i<�1R�o��'��Y�)��G����Ɣ��>�I�;���#���M��� ��l׿;s��4'(z�A��A �[AUE����;�.��:�x]!2h?���0�/�n
�!ĝ8��U�&�g����O�#�J6�yg�|dҷtb�KΠ`ZB��Au�ïM|G�tu��-�0Z�0R�l5)8��b�4؋���L�^oG(��~� b0�,�:L��"+;)�:�υHZE�ۓ�`ʫ~�;X����#V��>՜jf��_�ܩz߷q�>vj��`��p@c�.J���։�خwU��e)��/���l�P���y����dT������M��]�(��k�#�{�9i}ч�Po0홥I�cj�aW-�b������y:��Qq��Y�z}���1�|�R�"p���_3���U���2ב�Q8강��(����C�"�b��� ��P�?m�n� ����*1{P�s͔���S�9:�S09dqaH�ZT��z�2������$Ku.��*�J<�f�L�bAlmj}��n5c,�v�������[�6@�BW!�rУ����
~2��k��ۇG�[�~:�_ �R��6A��+�pdp�B�Ȝv�cs�S9��P�B�
����gX��7g�E�
\8�۴������W*,�Q5�
��rW��3�����G�m�x�`�G�w� �r��0��ʨh�Uz���D�����W_�@M^�[��)EhIZW.{��|(5+��u{�&��󓘊2�DU�m8n�	�� ���a:�`�8�u3g+;��ү��t��+|J��D�*�V�2������\?8�8������?3�T��!G��Â��C���& �IjP��N���*������L�(���[g ����8S4i�KYǸA%B�\�IE޾%^�V�W��:f�vݜ��)���q21*�y�J�~\R�F*�W&�Rj�}N3U�j[2���Vi��2Ӵ@��6�C�>�����R^��U�7I�l=�$V�x9[��4oF#�C�Q�>v�cQ�P���)���⬿h9߷>2��{?x�a���q�%�O q>�,��#���k7�*�l���/q��1�P��Ζ����>�y�ۈ��`A��wB�B�Sg�oE�+֓��q���F��:F��}��Y�غZ3��cq�l/��ʭ8z��[���]�r�
�ͱ�>I��X^�5콳�Y�,7�$`�C7W/r:n���f���C���b"	�j�t[���*�ۢ;��M��`���hԀ�C�d*�أ**�Z��/�5QI'���ouq�Xd��s}�����%�8e���]�#�J<���,8�E�D�1�٠'���v�e���]���?Nˮ�Q���V�1;����bT"[��Q�S/n|z�����O)MU�0d��P:B��͇b��w{Ct@n[���ݗ�J��)���	��^	��?M �9U�{:gl�����R�t�p@�����Xql�J�(b��L{��<�=��JӁD������z����*��D��7����L���p��,�`�(���ݸd<���Ο��\��� ���� !k��%�?���,����
�p�H ��x��\��"m�K&�8�v�<�DdJh��r�՗�f��U5'B��;���H#bfH��{_%� �KI�<K+��Q̸7wƀ ;>�7�
ʣʸ�/�FR�]+˼K'Q�.:�pk��+o���&�� ���U�����B�*�6�[ś�_4��_���`IVu_��ӌi8u�߉:�Fc��.f�i��"h�ޠ	������d]�v嚮�l��t�F�0J�Ysh�i& E����\�(3�R7�Ə2;5��yb��W��a�*W���өn1�C\f�r�k�`��!�����׼	�'���_��-��M�PP�������Vb�gC�tC1�m^�a��]+ɝv����6	}y/�S�sv!0�FZ�y�|���BXh`L���^��=���q��8'�*!
�E0w}��ssIot#��)W��9��a��30��� �U��g�\h�)u�du�b�6��uf]����р8:.�u��߽" D˔_{X�Sv�PTR"�d#PA(B��"q��D����qg�4�h ��_�P<��{�{yj��)�s�E�Әo`�Z�nE&�� �Na)��������uo��J3��d���@}�Ћ�R�����1.��1�nz1��L;�v��	�!�ā�2���6���R�����?̀�T^��ʢ݂4k���!ε'���,����n�aw:)��+���J�u�{SS��:�U_�K{�-!)Y<B�B>�aTO�uz6�;��<�U��狸���d��X~�^�X�W�7	ȕ_n��C���Hb"7\׹-���a����A��1T�@�9kCK4LD�������.׳ߙnu[M�6C��r�cl���~m��[���Qk���<jڀ�������'J|�1��Q����t0vy{�e�>��)�	/��Z��?5�R3�N�'��9b�uv��.7���l��
�}㠡����<���[�9����Z�(�,vJl
���0Q3�� ͚+Z��J|:��e��ɍ�~�il�p7į�:�:��g&՜�.Dϓ���i]iD��YCP�dsxl��b��)w���C����Z�\Lh�E�>���b��7&Zm[g]b����53�fO�x�C�kɆ)��X}f������BA����[��aP�o��{�d<�B���Q	G%l�9���{9֤ʆsG��ҩ:G4Nȝ=�Z�A!����|�6i�����
���r�Y�6X?���E$�BEy�b]6c@�M9Ě�W��;����"����l����y���*�ژ��뚐����������Ȋ���&�Q�`���Q�j	efY���X�[E	,!�t`|�l�6�H+��W�A�G�HQ#��X�.j�Z/�����<:�{��
��H�-sO��]c��I0���g�� }4���t&�_��K�9h�9Y&ڙ� �7>�t����fjj�=mx>���'��A�����׶(�w¦5	���b��<�ޖK#x��s�^H���F~1��:�n,�MN��[�q|��ar��4IG�*S��.}:����FR��)��
����f�iw�?U-�1 -����l�ק[�Vk&f��s9��Adk��g��x��7�����S�@*��J � ^���e-����d�nv�5�m��<Rh`��C"b��zWf'T-s}��@76��;UѸ��}H�tP>�}mP�_�;T9�0~^2���O����;%~7B~�p�0�x?F��r�w2N�5��?W�\�����u����$�
:y=@��t���!	�U�'���m����:��~dM�m�*�J�
��PzPw���+a�Fm�f�$�swʇ�*j�C���{]���{-�R|Q^�*u�lZ�2�Ń���������
E:��i	��ڶ���Ne�.��mR������� ���\��������˚�T+�켾�z�v3A[���A���i�D���)W��?��$��3�v���,O�m�]��>��w�g@���.�;�v B�RN�����u�q5�o�G*"��c�f�~w��]��i�P�³R3C/�܂����A��T��B��tH���'�a��4�u:}�������eG�X�kM%dxm�Wߛ`������T���.�����U�k�h�w�zI�8f�{p��g7����}����2�"c�ҟ���?���w�Fo�^]�ż�'�`.���%�6���\��(��^ԟ��Hkrm�K�H�VL���{y��֨C(9�='/{�Å~�RY��EF�K��lz�-@Z/$ Gk��E�c�i�|�c;�~�dz%t�V^���4V�n�P�,�h�d�A[!�`5�}���W�Z�ršd�ZN^���o�U�a��hB}�T9�v���cV׌G|�٩#ԛ~J	U�!��k�*���2��JC�FR�7b��"�ɋ�_�_9�k�%��U�'7����9�,#c�I�J3�i�����#5x-!)8�������G�x�
ϸG$�l����&�o'�	3����^f`�Jc���[^��ą	G�O�ճ���C�D^����t�;Ŵ9W��A��6�ū�Hg�"_L�"�y�7.}�ǡ�,��51#O^�h�YN�+�	k�qS㕔��~S����*��v�9�ڄ�ɞBl(���7���� �Ƅ+��9�Y����m�X>k��'=d@oZ��s/�t�o�k�$�XK��"���cM֗�J���֗�K�L�X�?.t#�W9@�.M���W3(�\S
��H���?-�f���8�>�B��x��[9-�����P��h����`-������y���]��g(4,
�\��'_�.I��2��KR�	� ���ކ��7}3r�B�.�L�q���"/n�0z��-X���B̘�bB����Ü��"\�������f�;�~ݩN�ƋtPz�@?O���$=ء�Kl+�@�M�j  D��+�� �R��7;�qX�;�ᬛ~��HwC��M�Z_��o��>|}�W^���=4��j���k��U�#������G�kn�g��ɐ����2I/{2�D3;�@jpЛ��M�L٦j�+{��f�ٓ!��0;�xI-o��&h$��E�ىJ0Q���Z�������l���2cq,_@�ѳA�d���2ʲ��g�Ϝ5�,C�֕Jݛ�WA�Q=C��w��[A�,�l��lr(��&�����8�]���T�2����x���"��-MN�����M��t�e �4�T}^(D�JPY\c���'��5E��*wK�pn���BYZhM�ڛ�Ļ��A�I1�kn�<WŬ�1�i+-��O�������ȃIZ�^�̝M��΍�^}��"q7jnb�D$��O����LFl�)ݚi��QGM��s�������%M�'��aYo�i����s�^<�L���q*^<i�Ӭ��6��@�(�l�H$�ޑ_�� �ƍfx��I�ԑhw+xM}��)���(z~n'�u��(��⺑;fd�r.�_�a����A��'X��f�)�=<6���3W�\�������֮ZsMC6�'���L��U����gI�����rJ�⨨.x�pג��HJM�KÆ���t�HT>��za�k3���&�	8v]��'����*d���hUvr�91iÑ����1h�4��cϛ�-2Z%s؈d,5�8�ÓbHP��������T���%�\��^���n�
��X4x�����Z}8`
��L^{�Dm��-���8��|�nCB�!��&R�2l�x��CS$�+�V�y�i�N��)6�9�R��7e�ρ���<8ؼu���Դgn��'�o�_�IM�ڒ�<qc���G-��m�K�\1�}��H�}}B��ti�xm�O 	�*�g;�S����_EvB���!��Ɔ$"f���
Xad!��ZŤ���'C�aXĪ�d��m#M����۪ʢ����B���Ш���u�b�(��w� �@�;j|��X	}|�.8cW?��K�:���~D�^24�&�������P�e����J�tY�g��-a�P)���jx�Ls�(�d�&1��h��_[UZ�o[5�X3�D�w!�Y����~T�7�����b�u��\����El��1Iv,��e)�ܱ�j�V�a�bY5"% ��.�I���a̲�u�:��<6��A�����t�����ױ���L-�#cZCk����M�D�x �Sr�����H���ν)%h�9E0�����V=���rn1�,;��A���th�~w�Fb�vbl��5����8s�S(�D)'|�e����%_��W�e��ᧃ5��xo�,Ou}~�e��5Q��,@����n|�zGq:1m�=G���I�SIX$F���ֹS)��)�����j������&�b��Q��}��J�X�񊁳���D�I#�M�!��4�����h����K����%�g��c��8�=��`�`Ʃ'U,�{���<��7ʿM[)|x��_��p�q��ft&��J�͉��l���W;`����÷<�y�$Sȝ�%N��� ��dLD�8D��.h�
a���/�ƕh�o1�p�lt"���~kkOj��-�,u_�:�ˏ�!#5:o���R��4�a��D	�5v낸����J,eV)�|�qF��z�͋���jU�lhD����<|����k���L�~Ԧ�՛����e���$���#�@G=�%`��_z�ܟ^�E��Ź���?��yxd�e���A��4>3z�6l8������ϺR�f��Su�
(uB�h�Wc��	�_�%����o�kW�̄���v����m22�6;�A�M�ٗ�e*G����B�]Lj�$$Tr�bٍ�t�0�tN�Il���;���׍Bֆ`껏a&�]��b
����03�E�7��!v4K�Yy�ￗ�Et����鮲C���9e�Ώg�a��o���[���3�nI���̃�� г�����et������sw������]�#u�Ԇ{'�{8�5�/��#�������d��#����{�f��� �x�\Q����d��l��H!�@����+�<@pv7�0@�=U��%�o����F{�p>���h��7}!.�wF����AcqK\� �)<�L�����.9�~)9��ޚ�Ёtl���.=�N��?W�KȆJL/�R�W���L�<�U�^�;0�����8�2+w}AN� ���Zwi3]�Y��7DI���Í;s�&��1m�هp|�2���g������Xù��FL���o<i��T)68�K�ST�i�Y�+��(��#����Q�6�	P��N�|�����Υ���Cj�1+-m_�A��^�wL���گ-^Ʒă�euV�,�T)�T,��-ԏ��E6�s�w[����m/�IX���L':뮢}E<�� ���4{�n0��T�5`=� ���ك�vi=�b_�-�~�U�m]^Y!��c�^�>�X���1��qV�i�[v�N� ���� �6���-X[�;jP&��@����,P[���Gk�+��#g������!��}������2ֻ�>q R��;��J�n�A�|f=U�\]�Yb�� ��������'�6
3�w�����Zp�\�������F���S�jU�E�]#,� �ӹ5��RX����D�äU<Ԑ6*3����4^��D�<;{�P� �������T�:Ģ���-8o���=oNv�NB-/0�x��R�g���s�p�ha�m ـN�����'�Lؠ��~�2�A������K>�ɒ����͘�h���U/n�P�Q�Ǽ@��U����|�S:N�]0����d�.��eK8A-�z3ཾ`p��1���o�������$q�0�[07m���4��ܿ{��>Q����s��͚ d��I�d�l�Y�
c�������E��kc(bI�5h��:d�:۞�v84�_� ���@w�x_u��EŎ#�0�jb�����c�Ѓb���/JQ ,0�+�Pܠ��w�1C�������4_9ad1�W3ed@�=E�_j��_,)A �D�,�p�����-�P�j+>ݳF��J� ���bV��B����z�W� �W�N�:�3�`����	��5u�x&:������ʏ!PP��`惡�/I�a�w�;�4gh���y��(�t�|Gj�����i��<�2j�b� �嚬�^�K�G�~y��^�K�l�A(��������/���?�*gJ���m�Z"�)�F��c%�N{s�v��dw���nqǅAQ[i7��m�����E����(��f�ډ9�92�8��~�j��c�M��dM_B��5B��Z���AHy���q�Y?�e�"�%o*
�^�v��<? �<���M��
�dB�U��3
wٻ�^���2@+W�f���Lq\K`@��g��B
�r���x�C
�Ƿ������#��>�����U#,��{�.6ǃ:�C�����UW��A*�+�	��ߦ�}��4��P]	�@��U���/!0����}G0�*{�z�nL|s7�`"[�P�T�-y~��,�!wˬ��|���e��Z�>E��[;��Z@q5RP�R�a"��ѳ�x>����Kl�Y�jG���F��$��B����y*%[���i�.VE`��`3S�����a���z�$4#�G�)�1ap�F����&�7g4;�c/�n�:BY�>l�tC�%�У{7��;l�e�|�є�I�)D�7
����ZF��N7�(xc�?���+����8����t?��������HW�ZU=�D�l?9�0�A; ;)�5�������Q=l@�K�Q�*v>,~�i҂=�4�s�WE!��C����C��W�~J��W�`��� C�'��ga�����9X;$ݮ�0[&b[�����4ٿ�K��PIB s��Ϛ�*N�c�;�q"?�� p)�7��f�-h��<�c����̴z���ӯ.V�WT'?K��<FSDB<+o"c�*��W�����⦥�R��N������{A����@v����3��\hn��5kˁ�&�ϐ:Ū�tG������V�Dk��w��х7�pE���d(1$kz��Rps��.�����~�E%W�@��֞G\�k����ȗ� (��4�>�I3d13��"v�� �DvNqI	1:�uׯP�����,í�����q����g�[3�na��B�Rߧz�T�0W�yj��u��7� �;�`�5�����L($��[ d��]D��+�hOO��f65z�V����f��<vD����0��\�<��%p��A2���*���-��(t��H��w��Z�r
@YA:H$��~;IC�
؋�
��DO��v{�\;�������u9Ψ<2E���~vY>����b���$�f��T_� ^FUSF^%�׿��L|>h�^����`o�c��XD�?h����<�p"v��m�1��?�4�U���Tw
��������N�7s/C�<
	�y{�k@����6���*��+�)�E6�)�����~�i��y#�Suc�A����#+F�@3R>�V���Vw3�t
�-���8[/ȅ�&L���xf^b ��O��^�J)��4�T�F���ɖrr�#������A���>&gM�#�%I�{f;��$E5���^0q�evƶ�A���'q��P��w�������ۂ_�'�U	��s����qr����:���M
K�f򺤊���>��s�m��2�Tn`J裳�Nֱ���+����*���Y�Z^�]?�A��_G�76.s�_�'�^ Q��1�J�e����z������Z¸��*�U7��@#M��aE�ǡ���}�G�Tr����0�$2~�8X��	=����Im�>�Ӭ�Ô'4�"��ɓ�����j�t�1��RU�HP�E�9�w����FH9�RP�c#=4��^DXT�0̀2����P��k��E�,1��]E�K�l�W�켽�B]�P�A��������y��>�j�,-�! ����=X'g��~Owi�߳c7�����%�֙VU`b�)x���2��Na�j���4������gp�qʪ_�ۖ&b+9���a�?+ڬfn$̓R�S_�Ё���rkՄ$8}�Gk�k�{}!yI�3�#{n��G`�����4� �cU�E���te�L��&\�b�� j�˅ ��b��zN7�ob!`�t�%_X�5�!B����b��ZT��:
$3���X�CGeᢵ!*��sSV�W�_tP6^�6}�����4Ջ�j�)j�x)�E�����fOi�-�[�F����B�gbg�`
��:���;Z�n�Xe���	��zA��D�Ff�fg�W���-�{*x����LLv���S{��?�ܖ�����ު�DJ�#B�w�(+b�5e�S�w��J[�VM�G��)t �?jo\�h��ֽ ��K_I4�t��7�_���������-2�=�H����la;�H�[����c���b���;����9�f~���G�I���]�X��t���ɍB�-�[N��;��M��!��:�ё'* ��v.3L�wEv^��z�	t�oE/ϼ	��i}���w��y�!C��=���p������2�^��/���~�˭ƕY8��J�Kt&L��N|�f�,_�"%d��(+:q%�A�%U�{:0��4-i:jv	��6/��	͘B�+�D�}<�_�?�=v���o�g.����m��chw���	K05Y~�g,�'<�>����4T���p�z~VT.e��<[2�b��#9qاq� ����7��ϵ����e@|����H(G$ǖ?�Y+~��I�椼��y���vNi�Jh�U�@��`qW�P�j�Ot�ñ�(�)rS���������&ȗ u��=ޣ��T8����w$J�'�,�JC3Y�gZ�.������q/�&��Uqyf����>���	�
���%�8 �����e�aO�W�?�蛬:-Q!R���qrl�ӵ����I�'#�9��x�,QCBy��AD���#���s�`Gf��$u��.����~&ED���!���qrI����A���$x�Z'���S�*�g�=�����V�ʄ�ZN�>vz�4��[��i�؍H7�*�c�O�a��3��lHv.+g����~<��{@�; �`�@2��g�UI����j����c"Q��m�r&0�?�	E�֗���ճ0��wߞ#��1�H�η���\��s;��&Ǖ�=�V�gH��͌�7
RP��ԑ�p���
-���m� �D`-iԏz2��Ø/r�f&Խ��迕�o���XS�1}-_��}��p����(T��o3��}�S��֘s�<wɋ�}b�("������y�Z+A}�B~F�3��d���k{NbOZċ����T\�6�:�V�(����t�6�\S^lƔ=��'�-I3��6}�#G>R��j� O$K{������07���H$Þ�,��c�߲�A��򻾟S��Ce���j�u^<��ٞ7��n��	�@3��jJ��A��ow��4���o� �@Vŝ?z�r���ȇ��_��O�ݐC�)��/5� l(1��잭��?�!����U6o�I+�p^� E��ysv7~C+_ёxFj����wDH9%c�K�x�jN.ق}b��I{Zp��y�}�z�1��	y��&~��SV�i�P+�G��o���nR��E�i��p@� �����T�+��k5G6f /8^K{Hi�3�]�؍u�X��S)WuZ�Ά;��<�����"�"���Q������8:��� ������#�M�oL2hZ�S�P���/��\#hg �,�q�Ru�I��_�a�ѱX����^ST�5z�����ac�頇�{�s/�J/��D��ӽ���rn'��� D!�K�6���/�XCc��5���g�:>�?	�:�*�c*�7W8���.�k��{���ˑ2��/z�M=���\��<��eB�uȠ~:�:A�ޞ�N{/b��������о.���ݾͳX5�1j�B��x3�Ƞ�pT�0�s�d!�R���nU����g��䮓[�j�׶+�#�G�4��[U<��y9ᨉ.TKQu��⒏���qt~�W�>�ah5K����0�U�s��yCQ[�<[h�}�_�h�'�w��/�9`o��w�0&�^��ͩ�=�[Q�p	���Z��}<ǃ�y��g=�ʭ�����HF�Pv%3�+���B��Y�e�D��JQR��Z�ջ�<2��P�֟?3����J9G��b�X.��F�g�"Tk�eb�o�]>�x�OB�׮����Kֆ�h��y5<h��No����C|�r0�If�D��T\�8�Ƿ5T���A�'ߵ+�A=����=D�s�м�bd��J��|�gI����G$/�>+�N}��� c7Lu��gz����)�!��'�t�v���莩b��o��0���'K,����\��5��^Y��.�^zL�Fl��*�vҜ��e����?]YN���q~���YN$��=#+P�e����������㝠ք7/|~uI�*��z�u���z �"�K�G�Y*�\���
�Y*�o�UN�y����d��QvS����jgM4�c�e�kX)�lGV�V��	�(�X͌���� �1���*�kE�P'"JJF��%"�#�H��(X���c"�l�$V.�10Ӳ�A��$�|�l��E�jk�C$0�~�@��/�Ӄ6�d�?�dɪ��v���%\g�I2���@˧��߮�&S?E�Z*!��z2:aM�͖@`��[���|�=��3+���mϏ�<t_'Oh�uwX�`r\v��*0<sc����?��� �h���춺{����A��V����I�/�%�{�e��1�圔�B�8��oq�
�����9�"<ę=���.q�K�loda=�Ϛ�:q,�U�n	M>���y��96�3��}��:�P�[H�;B�)$7Y��}��(�L<��D�Y�Z^������v�l��>�j �����n�9`�|�n(%-�����
	�J��d{�y�Ӛ����wE��9���~�C~�e�ti�t�Hyx_vXes�:�ot!]�/ER}�U����T��p1
(�m��';�+��i+X�x���9��kF�ve���f��<9�8�K60�λ�n���M��S�y\�E8�N�����?N��*�x�3��цlI!�i�괉uo ���C����M��W������rL��=c�4�4����np�`cǜ%QA��B��|��	C��
�@ڕ�묐�B�1��P)k`��w�T�R0�zN"�G^aϬ�n=٠��H#��VJ5q-0��j�_�8sx6 ��R��gc ?:.H)4Q�����
�y�hp<��+[d�Z�r�f�:_��E�Y�G��@���L���	|�'�5T�-��;Iyl~j���+�dCRO��3��o�|h!�2MN$�c��9-����+s��
���.��Q/SlI�����֝gk�+ݓ�4�>���YA�'�8�~kj���<�8���	�K�V�^!�}O^cX()�{
���B���(��1�ل�������5}���U08ә~���[WOl��߮���P<�cV�e
�s�-���V�P �1�l���Y������O��T/[�<����9�#����SVWH�ϴg
��ף��9IC
)�tLKj�~ueZ�����ԓ�	A��hO�{���W�P�Ѽ�@м�6�L'�P��tC7���Fɢ�+��J���ɟː��s��;O����o���
*�x���[埓j�:�I�t���}v�����h��L�6��KJ1�B�!�1���q1j�牿HY�о��+`� ��?�i����HM~cQ��&���Z<�UU��6�u�����Ջ��
.�-K��'��#��.�[��	����.B�e�ɭ��z�.���c�
�q4� 0�P�$���h;mA7�l]�Ñ��&����-f���g�W�e�;Dg� NE>m�1D�Q�F*I�ǡ��p=\�p	�|��~�g+~_�c��ȯ&�jwd|*^e֐3��2����$�a��0f��%�@��j'b�o㢠���8E���C��*�FV���md��tMm�P;�T��Uϗsm�1zyi���[�g�Rv�Z��(s���Z��y��yL�L�|W2D��Aˡ0`dx^��i
ͦs��h��v���2B�/�l�oA�o]�S��8��;zL���m���w����1#)��ON��Q�1�U��S/��ݩ��6�88�o.����:8M���"pdn����C��t4�P�P��}����sf��8n'ߌ(�Jܾ�z�'�,�ѰEi`��4W�*
���H�q��a�$�� ���*�"߮�;_�$c!�tܯ+��/^?�?�T��1S���5J:�02�֪�n�x�B#Y��j�3zR#rm���m����rٮ�}��y�����f�y�~��ɸվ�:�g\n-8�/��,��[���h�Y�>����W�Fr����{��R��E}L�y���km�,�b�%?�#��(_�O�%����O��:ӫB��߰���@Ah��۟����"b�C�T�4z) ��j{P,��5��[�V%��-��Ѱ�ki��-:�nZ7����l�l�.��fRL��g�I����?�bS���.��do�Nv��Y�c�\��<E7i����N� /)�)��M�6��SHI�d��6�I�f�fJ���F�J-u%x3�5���J��0/t����_d���r�2��e�M����3v�F�R���Q�G��;����Tz��^��[��un��~@I5�#jo�0败ڤ~�M���}����r�t0��f��6�&;E/:� �d��1���ݩ���1��wK"�Y���:S�(��0̈���'��͆�W2������l��zz��mV�a�C�D[����$Q�מ��P�@[J��O��΋H�L-?�h
W�T�����po�PM���?���{\ye&�G;�?Ag�U �}"^)���u0[���_V���m���)��/��bN�фmv�鏭�ڀI���^���5m�r���4s��P{s��3uf�4/ab��Wٶ��u��0���l��H�1���)�;������,���_�����w

H����<�K�� �Ұ�LEqc@|$fm����$J'z�[��k���17)�F���E�<t5�i��|���N#���KR&��ի��1_ Ћb ʼ�q�#���v�υ�S�	��J���
�b�ݯ�Y��M�}d�1Hp������W��"5�e�W�(!���@�@�`l��s�� pk0t��]�8]b<��@���PX�;�I��|�,~�z�yu��t)��h�,	+W��g��y&�T1*���,�qRl>�ؚd����5�F	GZƺa6���� ��M-G�h,���r�8����� �����AN|X]�����!Yp�Ȏ̵Y'��uYo�SUE�������|�/S��ae�ݙ�>��%�̕��.v�O.�9ܙ^�W0."Z��Z䬜�9�������0|aԥ��?g�"�:<�/�5{pRl��2C�x�����H�@e���%�)�K�i�d4\2����ӭ�'�ǰ0�|.�d��(c!��&1dĨ8�X�D��FɈ�B�T�K`��_��ӂ�L ņ �Yx�ף������_zSv�Ň��B������0#�AW8�..�s���N��z��/�^����sh��uػ�ٵ��!޼���o�Q�����.�:ĉ|�E�)o<����բF���i/��d��(n��~z�1�Jo����VD��Lk��U����}��<B-��b�.��1��iC�B�w0?u+�Cf�'�����cG|_X\Z}�Nޗ��+C
��`z�b����ݬ�6�$���L1e)o����流���PZ���̛C�4�pR�ɹ���RxiUv�c�U9�Q�Qc�;Ō�� �M
�s1��T��X�,#�&�cv`����Ay�͋�������?�aoa{����e��4��sX�S_fO-�3V�`D�ç����O��<A����7�[�Ύr#&n�gB�����[:�䉇�M*#���Z��v!����l�Rpj��Yȅ�J���g�̞0|�S��]g�|���>�"�)P���<�T-��7S�׆���3^0�]fI0wutRa��lvv�#�ɏn"�J�M��%�݁M8<W���a�j)���j�A�AU���u>�I�BΨ�:�5��~_MG��=��U/�	��䔕[,���K�Z@?e���&Ӛ��1�ex���/O`H��*��E\�ƽ���/�Z�hX|ro\{�ݽJ�th�c��&#�\����*hf6�����Nn����B�(=��h!)<�
s��ڌ�eY?�����d�N:��D.F�N���4z��:�����a�Iz�.`�s����LC\�q������:��hwҹ����P��:/)� E~_r�RZ�/������ԻKCq�{Qa�R'�ȀSÉ�^Nv�,��&�����I�x���!���o{Ha�Z\�q��N�l��^L�;���JZϯ� �	F͍������r���c�w/�Qu����<��E�ãmC=,����8��L����ab����.���h�?�����\��O,��n:R��y�T������q��	8G�ذv��2��ØA�ه�o��ug[�J�:h��"qv���e��Q�����D��p���}���#���c�W�C�%Pq�����L\'�͎��[��
X8��mq�x"C0k{���
�* ��C;�(3�k�%=G�_d8d,���O�#0��5!�]7����\#.�-�Y�ȌNٝ
�sϋ��D�r�r5����:ܮ�+���1��ę�Q<S{��(_��?��V��1V`8�	��E�Elð��Vu)���/0-�*�Zr%vX4#��[�^>"Q�p���j�,D�Z�	�p�70�:F���=rx��2���n�7-j��t�4}�]�o]�`܈���"of���=W\+b���X��A�賲h$^�q����D�o�_5+()���Lg�OQ��Yl�{x 1x��<�$FI?��ѳ�_��'eF�i�W�}��mv[�w��l��p+⮤��l��O��G�,���ܝ$AQTJ~h���H}!�|+�K��ĳ��:~�mtˉGk�JV����g'%ybC�H��)Od���-�&1N���X�ફ攵W��Od&킜*Dx�0���C7�\��T�9��C�`!�Ӭ�1��T�l��q+d�t�?�q��ӯ�,�.o��%	��;�}{ȫ��s�نɀ֢b���S0��'�=�g�J+^۷�|5�Hq,�s�$A��9�l�R���'U}�!Et�x��[�c��T�k�96�碬n�|�܅;��rQugrrQ��4"�͎}�c>E�߀j �Js�R��>)@�װ�Z6��E��k�f�D�� �b3� �X�M"M�h��Y��P�^�,W�6�e�vk�H%����:�9��ɥO�V�^�ך��ś��K�8.������m��� o��X -�Hm���&|0aϹ���L��ot��Y,��<<F��	z_�gB�i�����B�IS��k�g�{i��%X��h�C�+��Kp�̾t�Y�Á��{�C����y�W�7�m��x�鄠'�ܹ��EӘ e�<
�2��l�����]o��V�Ns�W)�I[�|�����$c؉�j�S�a��P��)?5�!r~(�p���_���	�n�!��sN�lm�V<mKl�]��Ix�Q5�3����������h��\QK4u�/�}��� )~B��&"��_���<�|�f�TD����7��Dk�ƓO2U	�P�ק�9>�w�S"+z&0wF;�c��F4����ս�}��к��<,*��-�V�m�Ԥp���5�L�i^�u����BS��S6��\]�[|��جZ6�wAI{�deJ�	���S�'^֧�V�(�8��d�v�F1=]�*,ul����(m��j��M�UY�5j�qE�cd���F��|�W5l *!2O�k�
KNq��Os��#��:	���91�fт�a3P�����`��Z����F�?���X�W���1m�~���p�(���3�1�6��YV���R����INƾ`��Д2�*������遶�G���AэR����|�x��-��K�'���m:a䈋0�֧�:��.�l/�^�iYv�^�m�{˨	S�sehB^��~;=![�r����h��]I����_ ���߇ۮ7�&�����+~��5��-���~js�� �wL�����$#��9� �Lʞ� Ii�|�Y+;[y �bS������1�Ĳʆ�=��l�>w����נ�>��aح�+j�Śv� �]�T+66�x�\:&½�=��,ÂI�H�Wv]^�ʎt��⽀�:Z�Lg䧫 g��g3D��=�&0�by�t�z��^Y�p*/a�r��9�2Q)����4 ���>�bG*s�Cӌ��F�����p�?hU��=X Z���c�,��Z�u9'T���1��A�%�s���܊}e�|�_6�сۓ-��Q��0-���A���&����gk��&Nu8{YK��R�f�n{T*�odc������͆_;^XO���Qv��������(�ue~Aٗ�P��{��P�S�?����(��U����9��U�;|�=F4��ö�s�Y,C�A�{krFM��'{8�;vp�k*��(BH�[l5O�=m Ot�eb�9���jڱ|��~���~-L_^���������on�A�Y����c}C��K��4+Ο��y=H����Bi��V`���~�S�E�q��DG�у`��R}�~�2�����j�-M�2nt0��p�q����Q�M��聬|;:��>�}���\;��1��˥\@��Y��z|�0��ִ��J����;R���[,�J���&e�C:�I� '��.����{@K�]��go~K�-]PϪ��ك 5��@G��m+ss�ɦ�_�;L�#J�%l���^������ �[ށ��� !f�_B�h4��b�C;3�Ki���;25�y�c�?��8�&>���X�������ָO��:"�����U��k�?��
rAW������.��+IW8�H%H�� W��_|�g�g�rzJf)X[3�Lφ�o7Л��E��C�_�O�����VUJz*󡁠O��A�V����Ǥ��ni�k�}MC75̊#����7�֝L$�G�������;	o�ըD;�.ܘ�����GD��¹Q��@�<99�3�T����N���C�q=�-G
��	O�uH"�o&�E ۷w����=*l/���ad����~c��5�ћ�ϓ�>$�<}�9G��Y���r5<D��s2�t����6��Yrg{�ᖼ�Xc7TzTXi
�g��a�?�P�،�0�-�H@w�T/��LD���N>�FmmY�������/A>�'/g;� QI���v�;^�,Q�Q	�x#t޼��ˑ��[Fߝ���4]𯬥����h�!+��.�4���d�)�������֠�ͳ�6�$n�v^���k��V�C��Bt�f8V2�P<��f�;���΄y/�U0�6���`V���*'x.2'�Q�౦W��Kr�QXmN7pr���B�ϑ�-�ScV7������F�/�S霼���ϋ5���^ğ���[�3).a�?΅���[�/$�K�~�fS�!K2��y�i]��vQJ ?q�}X��~��6�ۣqBa��+ׅ��"��.s����Л7Ả�	}���*�{Y���|H�
������ �7���c/��9%8I�����X�Ea��p��79�͔b=�o�qX�Z� ȋ�����~��-c��酡�$��9bSXQ�VNa��X/��U�L����QhV�b�`������M�U�ײø��׆괳$)kfVq�$ ��xSɋ���3�d��pKG����&)|_Q�r��Ӣ[�c ��͋�l�S1(79�{Y-�V��NG�wٽU=�h��oy3
aǲ"�q��|�yA�_��Amw
�8�Zk��9���ܗ�er���pn����u\bF_��n�0��Gg@m!'�$_͇za��1u�9�4�b��?���l5f���놋
x��
�	�F���\{w5e~�&�=���/w��=�ᚅ=��U^����M�anU�*+l2����w� W�$�qT��*�n(ZQ��d�O��T?�$��a�{��9�����p������Y�_�2#%w�����I�_lcM�+��R(��w-��Ɖ%��&�G6�P�]�j�sK\���b��D��z4���0_�%�%� ��ڶ�,J^OZG^{�!��'�2�&i.L�Q��G��3 ƈ�J0�],y��/:����lѥ�Y�R�V�"�M�X8'_'ż����}Z����cE��&�Rp�!�;�˻�Q`b�3���H���T� }�c�!�ؓ��Ď}��[\�&vv�Yd����P��3�ӑ�1��<9Y��)��o�c%h/S�� �A��J�߼F��"
ƍB�4�{�\f�jݨ3ibo&EJT��|UprH1���{�%�)�Z@�p�v�a{�#v36Ap�,j��8Z���o�O7�1?�|ra��I�ykcicoxa�����S2�Qa�-v2����*��Bp��9rO\CE�܍����~]Ҡ��.���(�f��Z����r�*�U�=���x3~'��&I|�z�Xdi�C[esd�|��Ox*�e>�������k��D��[}<y1G�!AZ{ p{x��e�"_�o�N�M�1� 'S��ڦ�%�D�D��Ӭ���Ys����7}<����l�Vz���d��#R�!���~>��	��a���ͤ�A�L/D ��:e�O|�� �М�d>��O�*� �����]����n'�3u>����P�ic�#���eu�[����8���t)߇��DysL�
YLp7<d�,[�E���l��Z�,Ϣ��W]a)�R��w�4�L��k�sH�db+��l��O)s(j��$'$z���Ƞf�Q�Wfݜ0sV��m�l���|�h@��s�AŰ�.w ���'�>���H-F9z��u}ɲ�q]�y�w����Ƙ[Y��+'v�����3X �ͱ4)̋��v�(٫d��|��z��(y��¿K���IyC�j�oi�c���˒���E��pm�X�q)�$*{�Lqˢ17w���6|�(ѹ0Y�Yu��c׽C2@Ҋ�KӡU
(�y��5�����%f�xS�ik�����^f'��� @<��:w���h��Y [v���S�F���:'���ɲ�����t�YAg]+�b�΂)_�<�O�Y�F�0�?=l�t5��!1�\W�9OT>B��(�l�7~tSFB��T���Ԭ�R-(~�m�D�O���͢%�����ۦ��ӹ��� 4χ'����u$��{b��*�J���U����A����������a����dWQ�$��{�#(Suin����gP�_�g�S��xc�Sz|�[]���G�=����/��)�ǟ��|v�2L��3������~-�V�['te��h��yְ�*y��N�M�ȿB�/HNQIX(<����T&m'f�޷���B��FIu,��.ˌ��(�k��(���Sk��W׊f�v��j^�8���r���k���VN�G -.x��O5�I��'��I����O��.y\s�·�ˬOOD���d4B���pٲ��
���9�L\x>��%��l���Й�6ϻü ����t�F�*�K��Q:*m[d3x>�;�,X�Pc�����1^��BM��]I HB��Ԅ ��2};� �,�p��i	%����u��+[�k�9X5���|s���p|z�4�,�����$\4�@Di6��d����Æ�����?��q�=�V�����s4bZ�|������ɒG�cMZB��f��44�'n8�.�i���sϺ��>[�ʪn��g;U����:�F��)�y(�ވ�p�4}�v1����/�m�٢�Yf�G[����I�����8sYT�`��eؑk������sE����t�խ��%u��8�3}�@,�O�������O&�8A���>�=o)����@�B��]�-�N/�a��۳I�*_1���L3 ��{mFܮ�oA�%�ԏ5���h�%��[��`k���|�Q�!|l�[�Wt�əL�Q�5�0S�7Ж�S�)|��_�HB^d�X�ʑ^�R&>�Ca��[���иfE�V��5&j%�Ǘˇ���롽mW��D?Z�7�+�ݟ�X��%m3H HR0nt�[�YHś�LD]>�i5�țD�s�����&�����o�|ZӘ�|;q��c������2cw�¿KU��6�vi1�����'��=o�����O㛇�4��i�e�R�H1ׇS�9�1n��h,�J-�!�*vR�7H�	i'8�8�ڀUa�(���Ȓ��l�΃���Y#�E��/2e*��:�f���ӣ���4��R��[����u.|�l���ż�ԥ��;�Ur�@?��˥\��Ut���;�K ȜGc�g�@�A���j�%㤨� ��Ni�3g�2�u�rH*���Pa6ߒ��:3�L��|��o���^,[����̰)����f0s�����F�����qց�W֦��&i\	DS�_�z/�~�f�m�ʉ�vfe�k�6�j4���9x�2O�Xţ�CT����dh��\RM4y���&�	s�<2�Et��>�@	�������vn�+�z?�U���'Bg�b35�Q^���*Wt=_ܠ	�{D��G�;�[�P�N���&0W�~,�/rˍ�[� ��D���#��QT~��$^T1@*-J{�S���3Q�R�t�4��u��0��K�����!Xգ���,�"s��������p0��:��MPCX��u��pe��>�IAV�m����#�M@�.�fd]�^�D#<���}߳<8���jFN̮[���c��~A��'W1(i0Z�C�sf{A��-צ���Բ�|L4kZ��It�����d��{�6�H14Wj+��0�Ň m=8(�u�ΆͺF�i����wj�	g�.���,�)՗Ԕ]��6���9Xv����&��T�o%��P����a�������_	�=zq�|X��A̴���Ԅ�i� Nʎ<�Q ���f+���8�Css ���ˣZ�[�i��%�jh�J���t�V�a�83h��oY�"��ش���Λ�m��`��ExV`w�pQ��*;\yKH�G0\%�	�u��;��s�2�$���I����6��H�\%(���K(�)�Ϲ��饬�%�!x�"�g�^ޞ�L�l�C�|&���
s!��?v[��/"ԍ�a9�����I����2���=��t6?��U,3z��Xy2#̿��C�v`�����??�@�Nd��K\r�K� QP�j�	���x�b1띙��.nj.	��b�"L5`�G���n�K���f훋�`\�fr���X��^�ѕ4)�Z\��%��/�Lo��):�n�����h	 )�$�V혆BgC�v{3+?^Lx���x�r���Y� )5���D�2�KMj���w��ǻKrf�ugAgE����Tg�>��-�>�t��ݙ�a�yܳ_w�w_����j��j�,�V�������c��&��"�F�S�V��Oʂ[�}j�bQ�T�h:u��<�ţ�#�I�c%�8�Q��C`/	�O��ź���W���
lZ^�da�d=P'�J�J{�|f�D�����W��|��H��7[����6����t�Ͷ�/��
i�0��m5qio���+d4��vJa~*��5.����j��K@�ݩ-�J�ŀg�Mă{�4�(�9���ǐ1⹙ڍ�9{��4~���9��V6` ���N=��U�sUX��ס�����+����V�Q�Q>J�!?�Ǹgj�<w�
Xǥ�Ȉ&k�����.X'k��\�w��؋���m��#i�A2�ߤ�s�Xv��}�fk h%���T�@����W~����x<B��T��k%b�w��~*uV��z-�����B�%^�茽�S4VX���A�ؔ%j��Hm�>��ށ���u������yRI\8�h�C�l�7u�+���Q�ǜ1�~��S�M�7Nq����s�t�2A��Ψ���)����
�%M��Δ���0]6��W/xn] �O7��[�)��bh��?V����_A�tƬd|���}��!��7����������kx�g��\`]f�.g���_`���D������z��Ї�3ă�:)����1�rDދ�Sbo�k0��z�i�=����l��ؐK�n�ZyjR���PPZ]������5�-��w2�P��6�БB��Tҋ*��j�iX�n���2����{��V_�Ĺ��)ad�wt�{��,��!KE�tDt��,'<<d�-o�t&����yp��zĠ�}Ҡ�s��*�}�/A�	������B�s�i 
Y����̇Ԋ�����1�ۻX��L���TBT���sw5(�͵6�Y�~sO.���B"wP���m�W;(����_�Б��`4�5�U��߼66�ҙr[߁���*�{�
��t:I�ի-�H�cs�"g&
�� C���LR[&u{o?n��8Y�=j���y��t���y���
�r{k21�G�E(�!�bhJ��^���%���!�����f��#�iuD��ݖ�n�n�EW^�ic�f卯���C��4���6s�%�g}5�3� ᯀ\�(Ή.��.�+6�5d'��7�����'ī�"4R����-栠>��-��c��9f�ǥ����LG�c�8��H��^�r�n�I�/�w��T��g��KN�4)v�BZ��*IG�I�e���p���+�ܘ���sQ�;p��l��x��XoeN��PE���4Sx�8�e�J�{N�H��S:����Ql�+���Xw? �'˦�Z��Ŵe��w�z���E�1��f��#z��a�[���s'nm�o�o�n���y1rԊ�C͑i���ӂR��x�q���o��;��Ug�XѶ|�	n� oNW�ڔ�FƍU:�-_�C�k�� zUˋc����n�iU]����P���,x����*"�?�-k��'��	+M�j��*{��`�_�ӕŅ%���,'0�)E�C�ƣ.Q�ޓ�\���`��֊X$p��f���H��'�^���xK���'�O�$5�2�s�́D�����m}�`��+u5Ћ�Ԫ������/�+/�u������:_�ߝ:��6-�lEh��D�������t���6�t�Vc�oW�&�P|�~-��x��y1�j�쒲�T��^W(I��;�S���gz_�� _����Oʍ��
��Q���5�_���S���$1	��p������A"�$u! ���ІC&�f�cm��e�6i	�����g#=���,!}1"M_n,�~���
0@[z������I���v�����lb��!�Jx,>y\_�[��@H�$���iM�d��Z����4FU������	R7g�BKr.i�'�6.݀�~A�X0���|�l���8X|��N�W�_��JF7�g�z��cHY*-�CV-.�6�a�����Õ��/³��c]����AV��
&���C�Zð'��3��(M2g�ρ��XmND�n���M0��z*St�'�I�T|�\�3����b��b�pqV�*C�*����}�5Zu�w|Eh���IDcJ�q���P�:?�p? (�~ȇc'�H��N��R7�붛CC�1�/�$���%�1�׍�US��P��E�|k�������1�0��#IM�n������'M����Hw���*y����n
��;��[?-����p�v�[3nO��܁��c��G�FN�]�m_�V&�BeIm�E�5�G��b�9I�a��0��y�ޢ���i~��P��D(�����v�*��G_�I�z7)�פN��k�3R$CR��+s<�(�*(��U�
�{���!1�`fPǥ�i������(*��s0�����_D�WV��"�Xf���w��o)c�a���Ls�Im���ի����R呷����c���ؘ��2��繍.A���$ �EH�n�e�4'�1]-��f�N�a�CAS��;�j%���W�n����`��Ni�7l�DJ]6d�?0�d���r��Kw���JQ8HX�}>�k(q��+3'��1"����əc����cS�B3d
�1�v1�W���+�-)3!�+1UXѿ�q �� �9����#�S��}��x�8Av�I�����"E�Hxh���8HG�
���Mg�u��u���))�<��a]Z!!pf��
G {�dp��V4����Õ���e@M.����%�])l,�c�t]�+g�H��Z_�w�M�g�Æ;����I4�	�x�� �	�'w�E�W6S�Z�=�0������55G���נ6f�_�g��rK��[,<D��Ǥ��F��I�7�����-8��>@����*t%ܨ��1��#�7m�k���"98k�
2i�E{�вs )�W�P���o-���|�e�r�"��ڗ��Y
M�ڵ�%����͕1�Ƨ?�KT�H�*u���j�K��x���IX��ᱨ�J��A?HR����_��C<�!}�H^���6�JrY$��ØU�aٟ?�,VRoc�т1���YS��3g4 '9�z���ݼ��4,%&�˨�4���B����ct���\5���:�Ȃi(�S
���I�nhX�ed���n���m�ٺ%ɴY���\@5�*S�e2�#~��ӆAa�50E3|�/l��-g��O3��*L�B��.ݟF���p@�&:���
j&3#��1C��|u�v�3��Ő�8E�a}���2�z�? �eHe��V�lQ]77�m��v.j��0t�حc��J"#�\�dO)�p��m2��y!Y�������L��%]�M�J4R��Q9%S�s�y��k��Uu"�����\*Y�e�U����n��%p�K3X~��la�uB�O~X�R�a2�aR�	i�����fG�1��#6���n~��&b9}�Be�3raX��C���{�,�<�O�)��z��A�d��-^���e?`���!-�{�[<��տ.�gM��{�wI�N�m�GZ�df�7�����<,7��/�=��[<������t3�<CP
�RzI5���8r�SIOs�s���g=묾����Qtp4��0�$��	ર#&�(�i�:ZӬ��ѣ:W�2�"s���4{i٩����B��_���U��H!pn��l���m��R�`�̑�b�eQ
{���G�d̟��q$ W��
��gVQ���BLBT��=`���jA�(�u��*��.WY�n5�!E?�:�*�vW��-�O妪��V���M��AC�c�jo���,l���4�ůds͹2p wTOx�3Y'���f��-A:�pqj��(Qω����WJa�uݹ�jz��@�/�,��tO���3i�:2}ܐꖈ�e���'i��y�i]o8똺z���+x1"n�>+#� �T-y��;B?#|�Ԁ��̉SP����T<�l�0�^l@z'dΧ�ZV��LB0�frt)�����,���1���g�dK�"u�Mv�ԏ�#�yq��Z��"�QǨ)�W�^ ��mR�{���ɗL�<h��]� ���䣋�t-|�-�_r�D�l�{�35�$�P�jM�������Dk(�p�?r�p�Yc���yD��Y��t�`&A?9�,Í}K�uq��	;$v���c�kN��?i|~Q�m'�f-�} }���K��8���	��֨(��
;�
����?�U�RE���M3������WS�w��vj� ��A��j�je+Y��9����ExFc����6v/@��������tT�����.ҧ�ݪà[��cu��V�N�7��	���ݺ�#
pY�02�N^z�o1��r)w���ǁ�U"���Ďc��G��5�|~UI���
������Ւi�����l��"�;��s����"G�0Խ��L-�h��6��א}�S�ع8"j@n-H}c)�� ��Џ{��,o��'y.�KS�]�R%�m~��҆��ڹ_/. 4H뾌B��7�D�V]�tN�+"��,T��r �!D ��?����2S"S�Ȧ9�Z���"=�t8�VH�6_j���g�D(��jJ��\���!���&B�sҗZ5u/	�u�ЅY��͕b�f�-hf�O����
f�͛1��k�=�2؞�A�/��K^���?s��bK����3,��z����XC��
��G��4���.Ӝ��˾�3a�(`�t+�nȍގ�E�����AB�D��
��狵��8��!9P���?��+��xJur��:_B����9U���{T�~?�X�2%y�2+\32ѵѷ�f����s�uL��d �'������"5t�W��0�1�!�dy�?3\��6O�9���� 5~J����Y}%�K�Sk�qkPM�6�ox7�v���`) G�&]��E�[�1�����#[y�(gN�U@��7���6�s�",Ŭ���ņ�J��@���߯�P"g��"�E�CI��ٳC�]�Q�Vq֔�7D�", ��y�R7��q��7�� ���HEe�h�?�1<\��Bb�`�O�18�#g�����iz�DMЭ��ȧ�T�*��E8����'ep.��B�wAD-�Ѝvj�w��}�*�􋸑��t�>��f��i��9����+��r�^A�,�����\h37�p�����A# �X�2�j�<��R���1�'8��nH�rk~͓�\�-V�;;@�ِ�jOK��H�4k<�N-\�+~��W(���r��x�Z }$@�B�%t ��jj�p�QA������Z�@�$��`�X׭w����b8����Kc�1�b����g�+qՔ@`�0�d��U/�f���+Oj�A<��n+ǦKҴU����6�\-�8����t��R��l���RÊ�>+ ~F�_�BV(e�G�c��Y@�8*��b��].�
}�F[��V<\�n0&`N���Y6"M,����;���C���xMz��.8��^�'��/�x��Iq2Ѱ�*NHk���%u��%�0Obc��+f��]��G��VńCN�z$���@̿�/v�D�j����btsYFgM��6|L�!6��*A��������$�zA�W�bF:\w��������#�cu0B�mC��W"QC�Z<1�#V��!��EwwELF�&\��uGܥ�D�?�Ior,+S��?u:n|Xd�M�@���4�΢[�������YB6F���P�:�K�OV�~���1��"�>�(p����U��=!�[�p"G��6a�蠇y���
}�0�ɪd��wTh��SF�����2�C�|nQ�:��`l��͕�G*���q�$;��}ڟ���H��̢�D�3:��@���-ƒ�4a�92��;�Ζ��?�i b�3�vk�M�3�K�cU�J���8�g�+}|��ǣ�?�H�g��5*`'�U���:w
�N��]��Q�Gy?��1�,|Y�C�XK7���
!�����ID��W�V�F^����a�r������`.&u��9>�!�c����E���U&ՠ����I��6&��,�Gh[��օ�d����j�1Wǝ�T:c����@o_**A���-��"���O�[7�P���q,���\TA�µ�	�'zի0�)�Oa���uS�2")�d{�GLl�K)`�%���o�I�A܂93�T?�_LA�ְ6T�x��b�9���f������*գ���gl���I#e�>f���iz�ǔ��C�$��FZw�S��C�|+_VhI�o���
\�-M��|��YwSg���������7����RG�$:��6��7DR�='�������I�1��������7��)x��dfi�GY�A�y.�v�:j�Ȍ���RA���iW/���y�x3H�2礗Zu*����).( ���	 @^:���9o�'[�ODB��(�Y���̷s�B��:.���S�.L���q�;�24�5g���l߻�_jzw��	��+���x3ho�i=�+�4}uZ�B83�1Y���&ej#��un�+ּF��m��Y���>��'Yt�tq�e��V��
�aF3�A-��r���b��H:��KDA�N�mI"+T��+�n�@Oƶ1~���O�;�D2x'�t�F�"=8��%f�X3	�0a�%S��\3�h������{
��<�Ђ��Ø�9�#��i������+���8�`f5�=�S�f�Yp��B�&��c4і*�ܒ/:���F��r9��=	��i�`e�ۛ:���O����^����IO�#����)�ڨΌ�kv�S��s4ow(n�@^�c���V���^(�X�U�����j���~Z��ŏz��ו��lj` ̝U��r�~4����X6qj[�A'�eԝ��?#�{A=@����P�gJ��:������Y,Yk�q���"�%ᝡ�U���/��K��YDh�s?�N45�t$���xP��ԣ��&�,���^n���Z������Ϸ��ݏK���?��׹گ�+���Ξx��*��5<��O�@k��D�\$c�#~,���r��`RA�Q�%�B�*8-�E���O#듫��ONQ��vH�|��di����^o]6�y0B6nN����w%�_��d�I�F	����i2j�~��A[�-{�"�1!�kc��+����F�Z��Ux) �-�Q_V6�M���0��^�^��7��W־I�l[�
����8kt/wQ*>cH9=�*%�.��QYڴ���/�b y֏'y�p8�t>�ċ?b�^�y�Ͷ��{�v�-���Q���6��DBX6˫#]Q�RθX��hA���X�uەŒ��@�o���P���oS�h�5��7�{ɒČg�⩔b�QH�v�ɏ-c��|���S�h���{��:&��s[/�U,i����Z��9�n�����_߈�}h�^��q�ں?�3|H|��~S����Tˊ�Ɩ"�bu) �)zD�cHFb��8����( ���<`�c��T�Eew�|4�c&y��q����ΧH�4 �� ��<7�J�~R��Ĝ~Z.������0<��y6�m���~�9���������r7CO��4ܣ�) �%nמs�y#6|w�m��,�^�v�@��^lO��U��/O71ȋ}f�(�5�Wm�Qt;�$�f�d�'�L���Mv����e����p1�1��O&vg,�����8_'8�4�|pBĦ$�'u�4��Bp�����8��>��:.��,_.��=k����ú�|�è>�ar0�ՃUqgLk�q�z^�"6q���(�|�;�}��4�\��ԳD��;�'Wu[�Ե��R��7<�M��ȍ'm�����{����>�N<E{ �9����)Z�	�
@1�va>IR�]���xѷ���fߨ���<�^��:�\D�%�ʝA�v��� r�8K��_w�z����S�Gk�]g�+6tnv˫�������l��7�Y��T�+�z)�ցR%0���Q��j�K�Y�J�"����F��з��JE�A{�TY�#Z�B�	��>t��f������w�/�k����i��Y�/�6�⼄|�(�.xd��}�$DiE΅<�T��
�;2VIbF�	���A�=?M�?��G
�tl�J9Zu\�Ro�D�����xr�y�^�ϳz�h��߲i�xd�_��&
�=
���w�%2�Al"�X��\jbyHz�?��?��)q��*����c��کc��laC\�h�%TT�h��[6*"b5޴!G%w�����iL6�X�ka"���-an4�lO��ba>�������K�d<dsU֒� ��*�%�WuҌ2ƥj�7�|�e�ɒd��E�	�;�i�	w_A�6�M�_��]��ͿȗT��J(��E�X��b9Ɩ���w�����Z����}=�=I���jvb�u��>l���o��lst*��YzH�xУ���김��� 0�*�Ҕ�5�ޕ05��Z[��5�pT�p�r��)�/���f�	��"�n"[?��R\���[)�^����3l Q��1�J}0<8�m{9�G���CT�h��A�jc{=����b��"|L�����v
t�2nT�Fy��:DCO���Y�0���ջ0U��0��+��ǃ��N�o��r�@�B�7�h�'	ɓ-�u��������}�X����;u�o����t�C�p��RIj�j�~E4/*�=�C� y�D�J�$���0���f�'>��JF�4�[u�qs�A���)Ҽ�F���kK�ٽ_�ciD#W8����f���pQPO�cVg����r��`�pr��}��/B?A�З7\v@!2�]yxSe���؉�@��x�{=�bA��۬ݛõf>%���h�r����G�&��j��.�i\��F� f����vS���%4b�	  ��i����#�"+I�iM�ه5��Z-���� ޔ5nO�Rނ�� F<aՇ!A�|�nؑG�	NA@N!ל�2;o�n��S9R��߅�7�\e�7^%��_�
UÙa龊��� '�|�/x~w���hD��,�c$.غ�s[�Z�s��g|�ׇ�gp(�7�����{��	�G��/(�����Ȅ+��a��9�{������MH�i� ���FF\n"��i�6]�M�7�njDO�4T���Mn�T��_�m�=�HO�Ni5n1D<�y��AX�GF�"%��J�n��=�ķ31��.P��B�����yE_{���c�r��$�F��:#~���gL�a������%��U*��^-����4�y�3t����b,��XH�wn}���J$�e�#�9�ϋ{ٝ�Oj?���<�b2�-* g�]1�wIc��%3\!��M��{1O/��|�=d�G-�L$!���8��SI!��ս
����ߋ;�qhb��.K߳�ep@@Ts $�V�#�}%N��X4B�6���%x�"G_Em��:t�{�e��e6��	z�S�3�d�ěy�E�jz�!�������`����Z�d5�,�8(���1F�\�'��jx��N�}W�����l�rv_�>Ё�1����$����(�,��
O�%r�BЖv��j8
l����H�
�.F�(���ݗD��Xo�V��8���>�4�w���RUO(��A�
����SO�X����<(�vѽ�������ֲ�,���S���1�P��Ѱ�+��E=�3_T?E R&<�9�#����&-O�#G���AL�Lir�(�������l;J�5>>N�8^�L_s����|JqQ�Va��f��fwV�ظ#�Dk.�Z�ۜ�����O8�+?18���e8�Z�#c�S�{�����SUnk��(�.ך#ȣ<~.y�c��i���̗�)�؛9�(�@&�s����I�ld]pqZHI�<e���ߞy/��߉�c�I�sB��N��b����Wdp�km��"R��5���%` 헉�՝r�TX'�9����3�Q� ��ū��PP�g� �˓36g�,���Wх��<��ۨ��Z��X��B��D[F�^
�;�����	��mi2�G����#�I��=1�,�O"�'�%'w��r9A_l���sL5	�*�3�!�y����k�Dx�C�U7K�:�j0K��<��Q����LZ�-��r�1+fV�Ֆ�q��v5*V}�_n��;�#o�w3j��mPv�!�3w��%W�hƐ_�kW����_b����<�bɎ��ӆ���������̥�}�"��;lܭ���t^:vF>qu��2Ҟ��Ϻ�(���j�տ*|D�4C7%	x}В
wP���Y�XOz����q$-4!A�f�c'J�FF�%�4�=�B�>H�������.����aib/N��Z>;�iU-����t<�z:,dk,.�-���Q�]X�����R���zX?����y��7�2�Ջ��-�غ���X�b�VǨ���c:�;0�eMQ��rv��0{(����m0�u��So�o�C=�w!���	�������/*����՛�ʽ��~��\k�$1;��X��hU`�!��3�D
� RE����O�]��Z_q���P�{47�{��9KO��E�V-�#��krBvhw3�v�t7��P�a4��(��ønΛ��U|�����c~hY[�n	2T�P��ѦW�PHGȿʉ㈡��{�Zv�w�����V���egO�,��ۊ���?�G��I�0�:������Y��TӯN��I�L��Z�}��A��CT��MAk��3��k��3�\V�<h틩�o7����,r󁑍Dw���H*�k�ъ {yx���Ƣ�W6tǳm��&��6���_JV�^�(K�&��1����+��*I�#J��D���i�ؽ`;��u�ҙ��e.��_��+�3���0t��0S���@�L;�K*v��8lۏ�鉚��{���ŔFTc�9̉_��_70���w�t.��p}��z���
+�8H���n�ϜT�|y%(��4H��<���|�!�/��*;��B��\LO��E��%���� u���S#=��>c�SR~��Pi.W����s@ߴm���>� ̪^z�B��{�a�ރ�˷y�v�ӆ�N=��#��$��1Wh�K�4��;�W�����ړږ7&v�DM_�4Ep������O�S3�[���i�E^-v9_&��2��4�lB��4F���f����,叭��N�/��1��e��0����c��E�RꚖ~��ۯv�s��T�ץ<��؟��#i������`��יن�+����UW��Ѣn�0/`�M0X%��>N6!:<�P�i3�쒛m$���p����%=S��g	�̅15m='�KF� �
�T�x��1P��e������<���8k��uTD�[g7���?
�n�*+�%��5m��a���Wz>,�`;Tנ�ř�*S#j��s0���=H�t��|U|E^cs9���>xV�����nB;?��o�/� lk�X�^./���d\��0oj��-��bvɕI:2ϴ�Iw��疲a"辰}���*�}-\��"o-�.�/1u���-�su\�sX�W����8��ki������Iƣa#q��)7��I5|�'���&���I��#��-`�#e?��������f�K.�X�2L����8���r%D����[Yާo��Z��kB�5+�T���JV�E��%�>�<.���E���y���D��K��F�����$Z((2�dw+x�=:��o�6J?б΂�g[	�PfHR���嬛ԇM׻�ܸ������r�=�6@����T^���>�8ZqS���BۍGK�`$�p�U&��j����'�h�j����C���1y̺�O�ڴ�����d˰��������xA�9��%�K>)]�1��)�5����ݞ ��T��ö��`4횼o��+f�6u=$�Ťil���H�7�y��w��K�%��K
d�����N�YꨂChm��M�&n����Tv��$&��X�+x��'�t���@�Ҫ����ׂAAup1T�V���Esn=W���cWSj<,~��/P���}��_c��r�Yahac�y)ɐ��uɁGi�Nd����KW#�'��O/t3nC ��*�	�҉��J�-�Bb�?��Mw��U�  �^����5���/�b���}���II~��M�ӄWC���ι��S����
S8��=O�����ȑp��!��������61m;�`��~W�/��ׁ�V�`�ԇ(���FS8��m���jN���5�����`��sz}r�7��y^��oS����y�w���`��Y�c92�����8VrsU��)�+�j���o�"7��8A5{ ��yC����A�qw�g�\$�'�1]KV����2k�����$�[�B(&&P�^OM��{:~y���� ^��@9� H��")|��U�h����D�;��5_��7�fs\�+�;���ļS�0����~2��.@?k��ڀ:��Xt�����F��!]C!��7��0�k�!�(�<��������KI���g�T�HX�#RІ��i9��s�A���ۜ��S�"�#�j�������y59��Ƕ���{\�N/��됇������<�8�<��^���~sbDIl�1d���ߛ���ՁQ]d���<m2�AcG����j�G/�(���	}��'��%���ȝ)w�o����Y�bɣ�C
L%fJ���}lY�v�Z$�n�\�]I��&��b *�-����eb��l�"cj#dl�� ,!�N�}� �	�~iP>���E�,Ʒ��3�k]�I��7�;l�y�:�wJ�R��+9���ϧ�/A���j!<�\�A�5�Lg\���B�+n�t2fB�{S (��cO�gR��kz�����s��:LEl�%1}��.�]���	)+B���4z4Ώ|]���Ӽɀү>�H��g�:@���OeDsׅ&V���-;�>��=i�gm��i)�@zR���51��uq������e]�y�* �;m>�vQ�`<C_�$.~�jO�!xL���V�Yv&�2��:���bQ�+���7��f��u������Jm�D	��o3@a�&7�bCy���N䍘������j�y}y�o�zk�z}��G��x[�P�q��-V`K���o�y>��N���Z��?f�S)?����fU��#D m?�1D�{ʝ����Oۄ��Ů}[�*�Z`'�"`�T0^	Opq?���J����F80�דL�_P�0�����^���
�ϵf~�~2�a�C�cG�ub��Ј���~���7Eg���Y�pb	��J����Ww�q
���DȐ;�����Z���T��]�n˾[~#y"�b;�uj:����x�kb��á����ߪ葃�!R�-\�r�D;��w��~���7��j
�:��@����w)�_v���x���L=�v�jl��iYƃ�j��p����wӾ����Q^Hj?��X�Y��[���Q�Z�
0��"I���(��J�Pߔ��z��.蘩��u�ҮW�n���gY��Q�4D X��ڛե��G�4���?�/t>ͬ�%�)"�y�k|gr�0�
 �>�X0���tR�@4	̀0���g��TM�ɇ��X��+�ƽ�t�i�VQ�wP��s�
(̮<�Y�)��4�$U���
σ K��=�v�Zu'�d���Ut����@��A����32�W��3�FW?/zݕ����@�)�WK��q�32�E�0=����4��l���v���0?�.G�d�%;G��� �DW�,	��� �V�{!��� �H~H
��f^r������8ի��zVΚ1�Fs���4$���a�Z�g����� �g���zТ���L�@�=v|�
�����b����4eC����:��a9:�;]�я�I�{czP*n����"��4S�vr��I�4�-N���ғ��Qҟ�4�v�+�<^�|�)�ȗ�=�C=|�03��l�����a�X$�V�`����;!��ސSc�H�~ml�l�䒲�����2�c've�Vb��
����5I��X��?�t��g���1�ԯ�
[����o0�Mq�T	ˀ���tՏp	iP��H"����>�F�%��[2*��1�m[�z�`�}+v�SKUBD�q�Ug�=;�<�s�Å���Ci�#n�B�%�w�>5>:�N���ZtUX��h��,�]h4z�݇�TT�23�|B[���]�:"�u�F`i!Z:}��w�=deI��L(����C܃�çz���a|��2�AfV(eiS7�gJ+���PVi�����7����`.q�tcG]Ad��n;! v*�O�CRMxе�6U�u�	�I��O�""y ��i{ZFt.���N��Io�N�?�m9+�T������έ�n8'^+В@=�,_��>�2}0s�?$cS>�-����}��F�zp����$��xrC��#��G9rͶ�搢��覯���G/�8cؿ:,6TD�2�ݑ!�oa;�TC�������K���%��.��@���`7Z U�-p��7W��7����M�����S�,?!�d��v��a�7�p�'>�:o������x0��*$� !�A@��'�U��g��ӢUje����՝�7�����˿W��c�A[]�!��+��ܭ)��F؝����[�`x������/�ɕ���zH<��2�Șj,�Y�$�&�ޢ�mqź˯�?������e��:S�2,3X/�EAj�)2tc��p��]�KT�.qm�T���6tFc�;�C�O�s�O#FXSDr����U���̂��z�~i͛+��j�gz�9Jg�.��l�����L��ji:��ت"��lv�ǃ�N�� �e��*bU
�mH/�b�Jm��������#��^�xV�L4�vq��䐫�����遛�ѩ.���qyX�f^@�[݇|�W�4��٢�?m�ڵc%h�1}�I/�0n��2�O����UV02_�G�)&l��dW-��3E�R�+>8DD��з���lNt�%TO�����,�݋�Uތ\�]�d���s.�"����!�b̪�5�A`��
�j	�*|�^�QͲ�q4�~�TY�J�M긳���@����QJb�n15����ڽN��m�e6c����������it�*4�Z=~5,�!�g���{m�8{�%t5��np�!�� +�`ל�:�CH��So)U��*�c(����B]�y�BC��P��kksF����9��V}/L����c��v��x����l8��w#
˫�0~i�=s�����Q��P�H�@=�{�to!���I$�b����A�B���y��/����hKc�%��&Ύi��>�8�d28��m��r��|
<�(B�)w���٨%�*��z�;b�'c}G�[�3ў��u��Ǉ	�'j���r��Ν������Ln� ��u�б�K�] ���Q�����{^M�[@�E�*P���S~��*(!��Y��̘��o�?�E����L%��ȓRL���˄N�",����-񕺤P'N�AQS�de����ϫ�Ț�]1�[�oh��M{����L]�"4j_�5e#qHL���+Y�/e咸0�fbkH-����_Z�����I8��C�;��xA�;��$&'�� ���@k>&~�A�U�����l�௚?0�	@t����;�^��u�u�a�1�Z���28�0����>��\���������_�UN䉍�	P�S̒%"$=�%�T�b��s�V�zŶ��8�����XY	��LPcgk��� ��J��kl��R雘u�"p�&��EX4�3���v<ﵼ�M�j�
�u�Ê��׬�!�vf��ؾ�r:\k�m�E띏l��p���(�����~�hɖⱭ��b���𹮱%��<�}�T�y���9ܙÒ��i�[}�^EN�!?��#�R,�E�3�\�%�џSF�P5f�4*�����C����t����
�;�?��d<�[5I�\c�-Z(袚��f�)�Z�4���U��
Wⅷ	�ܦ�lǃ���:ěFc��I�yN��7�I�U��CEΫ�!E3��Ü�����t�Js�D��f	���5negEP] ݎ�l�����?7���O�[��e6�Ojq*��*���l�-A��{�	!�b�����a�����6�gUW�V��-��i��� ��FK���?B��jh������,���G��v5c���;bX�?�ɸ�O�"5������,�����j�P�૒�����]�c;_�Z�l�I��IWĚ���u�`m�f&�S_��Xw7��8���N�C�/���$�j4���NҬ*���Z>_�+�w�.>!㚌�7���whzO�b�����8���@Z����(1���A�����b�
��352���OI����>��	��������N�lȫ�ʰ*V��tP���x3ޑ擞��` 4���qC&�i�G7*��k�渥���˫NZUx.�]D��n����1��I�q�\�
��f�u#�s@�kI{�7��L����(��htmKj$C����A���WՋ��O�4�;N���M�l�f�%;f�bI�W��	�I�6xR�?�I�h���t�����r��d���=���ѫ�#0?�(h�4�t�_�g,0�&z�ia�E	
��+�}��+yRY��~}��]
�#�~=��õ��ݼx[�D�C.�֧pwZ֝��Z�޻(��w��r:ƫ�,�M��S"��`�"8~��Ү�4{�:Z���b�����*$��#��r8J�о�k!)�85$�+��}��jM��2��5��f((�>��6N����'lB.�Z8O&��R�i�}jsH��bS��7��хUJ��ł��'����d_�PY��"-ߪl���w8�T���<��^�u!�aʘN%���f�9�#P=��k��sY��A�tY�KK����Pv+=�_	�5��}3�O�
okma���v��b����a�۔��*7��n��/˔�_x~Vv�LR�rP��vWz@5x��v]dA��Pu��s�	S
�u��[��Ț8V�K�'�a:�D����,se/�>���mM1������XF��K,ʮho��u� �A�� � �������F��d��j8I=v[){�������2+J��u�Y��Q��u�*��M)����@l'��m���T�c(-�YG�R�y}M��Z	_�<b,��ät�J{���D; I9�X����3`9n?�l�U@M6Bc#U��8��<��'s�Y��$l?MH��`��:.�	�<���`�]!���k������J76�F8�y�e*<㇡�.���䕡S��ǿ�F�h��V��#��~:+����:+�d�*q�Th*t�槷|+�v�E~ƞ�lԃK���D�/&��qfҼm5}���R/Λ��^���*}ԳJA�l�N���b� -Kt�1����b��0���P�]n��7��T�����RM�v�+�/A��]Q�P.��3���2xz�Y��u��\�r��{�w�w�~����p�<�|m>���!a՟_R7��f;���;K����� ���S����ΞВ�y��ԒvA�$W�6��6�CM3 ��j�\|DA�P�q���H��\{���|��[噵�x��\�T#��(vq�TB����z���{����yd�Ȣ�I��;�x��ih��SW�^���%���Q��t#e�=1�pm	;h����
6�'�,z�7�̑���շ#��(D4��<�a�����M���9k|T^o&}p1q+N�6�M����c�{�?FE�����C��J_Ay�Z$�3"�xQ�3�v�ԈcHk�w$�5�ѫP������q�����$����"]�a�L76�D4#�
(XIh�9��2�����b�@*��͵�_�2;���������*n�*�8U���)\/���@��jf	���xI����a�f4|�����y�?�A�)6���ϋz}��Yx]��$O�����{�~��IϏ��)��6��g~E��a��sD�:p�6�a�QJ��D#�`ls'�c���M+��c畘c��X,'y���̡mɺ��Z�U�x<������W�mQ��$��ޞ_�k7�ů�����i1KD䈯�`�h����4 n�w����	���b�7��}V�E��\�J�NLzr�j�j|ΐ}���c�W�5i����Y��`y�w���7�N�9mgL,a�a����[2�Q���ўƾ�F2im����V��j�'5���$���:I_��K9�I��/{3��W4^���Ɠnp��N�t���v�U[ ,��j����N
M�kR�Uo��s��`/����8�ꃩ10�&�F���B�^n�O4�"%0������Q�n�uuO��/w��X��Xw{s��߂U��Rue��9y&��1�.���{"�y�'�"
Qj.[2�}Y�|_�qȉ#�2sx���X��$lZ����pF�}h�
L��=�s��XM=�PW���`�U#�fe�d��p�b&��Y'L`���~|���醧�R_����A�`�Ҿ��4p D�1J-�i�ʫ�E����F�e4�u<:��E�d�=9�-'r�� ������Kک:�S�A��R���d;0Ww�K=�9��A������\ߕ���~�~J����,|>�7G_��B��1#-�X�kG腐�a�az/\��²y�H�(�QZ%&l��XAܙ.i�b��8�(�t,�%�d��5c�b�����G�b�@՘���y�����7⑵%F�u/���4��oZ3S����v#C�x�<C�3�d����c&"��.�.�ԍ?������o6�9�F@�2���G�����JxpF� �z���W>�y�I��{]v�w$[@�ʪ=h�����L�ި��`��Cԑ�D3h|�g�#�zEI�17	�k�Bܞ�"a2pa�/��j�"`ȌǊ����HT�.���B[���5P7������d�#�-
v��j6�!ִ�I_�蓆-�ZCo�7��tpC�c%-�� w����,ʶ%�#cj�̽{]J�Ţ�ٟ$��r�9�գwި�=q�i~ޒ�#��|`�����iL}r�J4�,A�]Q�v��bb
f���4�Z�5%@�J�R�����>��7��o��@�!9u1{f��++����_��~+MN�Z)�P>��3��3��"/	�#���4`����u\}��A�k��)���|�G2����1]_ y�	�3���@R4۪��=��o�� �Flʿ�����?��
f�(�����l����`�pj9^���������~{�~"��=��+��:ɏ�[�����t6����8Ɛ�����qȡ�����S���n�jS�xu�b01􏵨s�Z�M�c�ʚ�CP]Tc���]�æ�ɘް�7oQr�7\���"�x\
B��y��N�u?�'�S�U������~��ѭ����j��c2E�9j�;pA�}Ex[4e� �!Ď{��/t�(ns��<T�W��fV^�'��[�.qKs��[RL��NA5^�Ȫm���oAqXM��CO;�s)$t.�ሇ:�x�~hʤtL�0m�d�/1������&ƾA[V�@Ǵ�ؘ�e�e6Ψ�)m*u�W����h3zL����>,�����79,��0������ӈ��ܼ�F$h3��
}�X:�	`��PB� W@�8�ɣ�ޞ=����p��4̩5�M���;�7��+ɘ��B�Z������1*�U�H'��q��\?Xɒ�*D)�����aQ4^����\����~�ZzgM>��v�qy 7m�uh�$Y�:�~�K}��{�kj�B� *�]{�������#��3�A��kVT��zb��}��I�0�ɯnQ*��P2�����p�-0��"�S��������:��Z&.����<� ��_�X@�l�y�Х�Q?�ް�q�����t]�5���H�p�ʹ��il+O�	��	o���&���k��k�Ƀ:�8q��;:�t^9��R!�$-l(�K�
��'�{�V//ă+JE�i���#6i����oA�OIkŲ}����R���v��R����HPbx!b�2�R4 ����b+\ ���p<L�fN7e��쀜��#?c�G�P�>���	��&� F��_נ/g���x�]�<F����i7-�~�顮��q��?�f
��,�1����N�J[#���*iv�ӝ����XH���I�'&�v�j��?e<��
]5�xZ)��;SK��ĺ!+�zTn{�V�?�V��V>K�h�!�y3>�t���R�R���֮s:�z��n�9�Ԏ���j3h#��G�׫[K�kԃX5$�c\+���ˌP��:Ν����N��Q�뽗������):>��;z�2z�#��{!���`�x���U@��7��������������^��<�f�5.���Eq��+�ʝ5�Pi`[u1����>�B2ـ8�u<��%��?8 
��N[/ȕ|�/�6�*����E]ޖ����X��3�8H���UåVz�ʳ��&�Aڱt:M�,t�֜Z�h��.�Ż[����$:�jIe����q�D��Nh�ԣ�PԼEڑ����)Լ����QI�]@��P�����TQ�������J��8\;HO��#���Y��w������S�R�
������J.��Z�;��gL��G:m\�e��gtL�!��]�X�R.�%w�m���/ֶ&'mu�-�����O�ԖP3���5w����<��D�f�,��-��ﬔ��s��f�ie'6!�A�i���O([-F��Tk���N�y�3 ���aV��˃ӟ�s��iIb�G[5�D�+�ď�T1[�����uޓO�El�dx7B`�G�M�v����員���'�[0}$�v��,�H� ���͵���a�i�#�iuy]� ����v�jl?X䍂���b���*e'8 ��m�?�z0J"O�'�?e��s��k]���1LR��U�?�e�(؋}�6�.,`�v�����<��o��ʩ����S{����i��U��1g���H�#�������d����h|!{G��Q۝��rF؊��Ǔ�~Xx��T��%k��(�_#�zY��m��Q�O]�nB�[���K��x3�ہ��ywr�N[_��U�x}B�K��x>�3&Z8�I��Y�������l��-qm2��n���0b��b�Syx�xp��ln?���p�=@��UNA]�~�-��z=P@�_�������9E��FR��ޮ�� �&-�?=���ɽ�������������I�<�6$�Ŕ|��Β4I��8��s��+�m��ή��X���1P��K;l���E���V���Q	�o��L�%��q�p�^�A���OP���{\���������@�C~��9Fb^�R�H����cM�Z 1.���MQ��Tk}�C��"F:O�#~��7<���M'=�����)��؁<'[���z���
��+?�=N`��|e}R����>!5>�#�K}�Ʃ:/+̫gM�RŁ��-;�:�+S<o�p���X�Ů�G�gؿ��Eja�#�K/�N�xJ�)K	����!w����m���Q����&n�����H�6}L���-�5�7��Z�t~Ӳ	��Ep51>�l����a�&*�f�Q��SE�]U$�)�C�b?����o�H�D�E�h�}�6J/��/�4�*u��c��F;�_7�K���/@\w�;�z�# �7Ё�
)yW���A�$V$%Lȃ���S�E��8��[Y��a?�"�[�2l�Kg�(a�.��2Q�RG�j���ٺ��6
�'%�w<�q|��+�	A��F�kS�o$���\�.�I��Լg�Z��^�{�q�}�R����K?�<����*��]]������U3��	aq�|�/U�ϥ$��{���%2��K-MȘY3�S�=|�o�F��X΃�׮���!b7S�����##��t��<f��7~ܻ�`��,�:?f�W���buH�ग़�-���X��o>4�:)I���fM��@'�TS�6C=��a�v����H&,ހn�f|6F�o�k�S
F�bՎ�����Đ�q����O^��wԹ���>ԱĻ��LW�����Y�G��˿[�H�e#�����Ȑ� �j}ӼW� �2t~��I}B��c����Q�
\P8�M��b4a��v�?n������w_e��$��R�7$�l&sI�9l�/-8?����%� �<ؖ�R��3Q�f[�=C,��2��䫙1�#Z֙s�7����Ω��Ǚ� ����b����M�?�L�=�YUlv6�� 2E��0ڔt���-�M��wZ,Ȳ"�����Z�c�WVmJ,>i�k14rE�8�j�c��l"�m����CAɫ�4��-�R�����	Bͺt�i��wOm��pC2�mx�?�T��:צ<�ńCa��x¿3�����=���Ou����CE-X�d����
S�Ė$zC�abV!Cg�)X_R�J��}��_R�T=�q�PB���M�k@���y��a�}}|�%��G����H,4y���f�5��Q_>~@�3��u�B/ܚ�N*���w/A\K�u�����_L���V#�`�C6�{D��ů�.Z�!�#�!� y��M)ؓ��%�����&nJN6��w40֐�v�)+�"��]d�S�&�F.�6��a\��/�_�yL��ɯ�[Ѫ,u�m�R5�xA1�6���57�Q;��gܐ�al5z֢�\�J��2��	�����[o�4��QU=��5�\|�ʝ��G�5Wl�-�*��NO4�T��8������Q�_�)9���%��c*�o��2j�%��*�AE�ݴK�r�{'�����+4����l��h������ �)���$�n�..��W����9	�B�����>*��`�y��>����=�{�E�M���Bcd�LS�$�{ؑ�$t���5^z��C�LNJ!G�_���Rw�h���q�f֐ۦ�l.$x�� 8@�DiGҵ ?��r��9{
�.up������T����m���T�sÛ�8�`�0�9�_��W#s��_ԋY:F�����}�$�ޜv�չ%�,>��d��-;���W�r�y�RpM�CE�)@�b R�c�Ɖ8�M��\"��y�&\7���1�8o>O>�2�Pa�����S���)��Xg�U��!��[:�ܙ?3^�	��EuٸIM&� ���'���&v6�LC�1%C;07�e���v���&��b!*]?'����p���.=�Iu�t���!N�遜HB�:G�B:lB]�x�,�ﱾ\�II6d5����Ԥ_�H������L�l�Jm&�k��g��,�u�5�M(`Z2�L��1�`f�ݗl���}~>����������6(F��i�7@|u�:R�5�*9�u���8Y��S���l�W`D��������bۑ͕�|gW�2ݿ�'��L��6��?���Bw���-�Tى�t��,n����1|�	z(�D&-����h�a�7��?a�s3��%:���!A(��ZJB���؋�o6r�%ʂ���!��?�$0A�!ޞĒA���v����d�ml΃U�" �҅՚rz�I#�
UWc2j(	�4�,�����Wd1Q��u�*�*�=MU�s�.�'�9%�`מn�P􈠜,��6K�j�Ǖ �B.�@�)�/V��j�
����.!�?4���<C.�o�m|0�-�Ӿ�H��N{����ǵA?&�˭z�FH[�Vb���0�ტ����/�t��"��)^�o%��(��������f� \F��O�H�P*"�J��z�	4��,+Q�
�w�@��UL���8��8g��p��$����Bkڑ_3��S/��oZ0��Y�q��F�`�H��`�E�0�����5jn��
�ب�;�����Hw��@?2���1[լ�V����<���c�VbD]��H��<�ri,��e�ԮDV��n�(�b����r�X���x������{�S��� ��<u��=���Z�Ty<���c>�Л�@m@�����&�1��n�낭��wt|�`��ʶȍ���Z�D�5J �&˞�#|��yB���b������-�n���#]a9��ܻ�����J@�I���E�Ǖ��_z��F'��A7 ��n����Su~�d�͇Y�����=���j9{B&�VKN��`���z"�C�Z�!w#�Ndc0�����0>�=�_ؒzUK�=�J�t��"�g,Z��.7��m�_R�!}4d�w6r����K�,?���nx��h��ԕ3���JG5�B!��#�<(��e>�m��r֚�cc���w�V�7��2?�������f��88�`�N���4_�P5���Ů�خi���#�zب�ɊEB
̼�\ 1\���%�B��OҜu�2A��H��9b��c=��VL���v8��5x�[3���?I�e���j��wE`��fR}���MM���*t��h8��qtLb�U�$fy��3 <�i�s���33�o�llSGг�G6�Ry�$�(�??;*tb��Z���gou��J�A����T�{�R{�h'_g!����~�ig'�&@�ҖQ���V��q2N_�;����`�V�+u�H�D֓����o�)�)7��nDv�R��s���j!񟫘����j�3�7�ぅkߞ����4u,� �뾠�b}��O�٣���9^>W��G�B�ǜ��~�[~��M�n뜡����B/m�kn�,g����g�̔JN2���堨���� Y�E�a�=��ʝ�x����<�$=����V��(wL�����/���
�e��j�����x��R�(>���_$\�=PՍ��.N��&)�v� �c�qԒ�c�;�#u��TyeJWX��Z���A�w#tA�o�'ΧUT�?̤ޫ�n���	;��M�"��ͣ�K$@9����>�g�J����DB�����s�C�Ht��5�%� 4��崏*(���3E?V!�1G�����^�����h$!�J:	K��?0����}N�����q�p4����N�K�:#l�����E������53z�4�ᔧ�v���QA����5�`��/�m�����C��m9�iB�zi��+:~A�#��wR1��8�j�6�Z�Xl��6�p�} �)�5�"P~RZ�v�h�躷��_ƣ��ct#���y�$���.+���x���c)T����Lφ[�~m�8�F�6s���e��u�N�¬��e"~�g�ä���H�pnLe��x��g���ǘV?y���nF�Zҍ�Wu���Vh-��1t�4E
��3�c���ΰ)�#\G���|��_Y���X�⹾��Թ!��u�H������V�n]L�6���延��6�Ol�U���tvn
:��L�����8����M�
��'_��=lɦ8	��%ټP��K�T�K�dX:�en� 2��j'��� 0F��ō�ef�%_`o�k���'�t�xO~��)�.^F�Z��'眛�ʯ��$<k�\X/��H���4��?�Q&P�����$�<!ܝ,iq�ԅ��L���]3d���?Wo{�Y���^9%�����ԑ��Go� ��e�r�G��>ʔ����՞�Bm�_b,���8xA�nI���'�耂7���\x�����Z4E����n'�K�7Z���,��2-�
jMB4d�צ�Eg��gA�Y��+�&�M�w�"gNΎߺ	Z��V1J ��Z�d{D�X���C�P跠�4��>u"Y_�����n�r�/�17���=ׂG`q<V�l3���&+;���q�ѹ��0de�Dv)x�U���u�$T�k�Vحy��,�����>�tYK�?��@� }CL~�C����a{J �$q%�&!�c����E>ۥ�A�Q� ��	��%�W�[b�ƳFG�p�P�M��p
�����?,��vFQ�ˀ\���\�=�)p�����@����ǚE�~(�!Jfj�N3��{B1=Q�s2槈�D4eu1����+S�#���ͮ.Զy�W*�O���Z����k�ϛiG��0Qo2�b���I�e/U/��ܮד�,�6�����9t3����6v>��mx�u�7X&됕s?jL��*߻��>��4	j,DjkwՄ^kNf,mg���=��u��b:�$��y>�1���	��HO��L��>Ď����ƴ��W�)K�Ӟ9�n��Pa�C�s,�G��ϻ���2,�Om|�N0>ӋTٱn�l�@E��Xm�� �c����^!-r� ��p�U:xk��)^�t�]E�~M1�ԅU}�IzY�����͟�ǈ �;=��Y��:+��Iw��3Elo<ܾ+=!mTgI=��-R`=��9�r/k�x�R�c"����C�����R�_�-�M�fZ3�i����m.��6��L^�o3�7;�3�[=��+6Z��L�2�;R���h�d�.�ũ��?�pB�����vR�E�)�vs�Mƴ�ѫP�]��̪�����k0A�l�9��K}�$d7�o���L_���W�q4��ƀ����_I�}1�|O�FnIpxe�1� m��ZJ�ݚ7/LB`�֜kf.�>��
LlV�RF���~lf�D�������w :���E/e��t9ە� ����`vk����l�5��1���ZB�~����W;��:�G��u���?b��u���ͧ�eZ�K��Y@ŽTx?蟿,!�5u_࣎��}϶FM��Bri3h!kGX�@|���>�(�O2����O�����N�@���T��JoZ���3>� r*~Z0ta9k:��>�.Ū$,&�֧Љ�j�Y"�yso� �@���V6��C�=����q�w���-���	�S#2�"�>�fó��;T����TbsajdЍs.޾��Pp�x�{����Q��H7��:e��aG�7+#�Ң6>�kR��</6��r|ѐhׅW`L�G��m��FŠ��]����Xpe���k���T�0A�#Q:;���Wʽ�|�z�����JZ�M���m? #��崥Ԃ���\�,;����=M�=�LA��D=����9�xl�"2��ںdx��G�d+F� Q[��=ȃos-[۠����QDt�`��34�WZ�9��mr���̦�?��Dz��B`�/�s�a}t�p�>ΰ��f��G����i�pt���*$�k�vP�	6b��v�iRf�kP�af��v.^�}Rp��;j��!S!"w�-Y�v+��rޑA�x�U^�}�S�o"N�B���Ƌ��nT샩�H�{wjؑ�ZlQu8�ܯv/W�&��X�)T��4��A��Q@�u'��
z2r��çô�b��߱�8m/Z�ⶡV�O���_�X�H��o?�����ۗ�n�m�[�<�*󏁨x~�f����4?�U�ڔ�g�.�U7���Xa��N�oTv�<��K�^�����Y�\m�b�+).ꫲ?t})��3�����}�x�uS(_;��y�O7��_���e%P���γ��]�m
\�PJn�b��%80c��f>�,O�b7@���!1�n�P�r��4a|��N���rc�k�)I!�Yz~��F,T_rw-U*�V&�p�j��{�o�ti�'�ք���~_Ĕ=~�B����(l��f#C���Q*�x�w~��B���I�:9��O�6�'68U��'岼��E�� �"[�OeߘGb�E|,�g]|B�	ȏ�٠rYr����vS�����m��$��Oy⋈���w�X�B�!��