// cycloneIII_3c25_niosII_standard_sopc.v

// Generated using ACDS version 12.1 177 at 2012.12.05.21:45:54

`timescale 1 ps / 1 ps
module cycloneIII_3c25_niosII_standard_sopc (
		input  wire        reset_n,                              //                         clk_clk_in_reset.reset_n
		output wire        local_refresh_ack_from_the_ddr_sdram, //            ddr_sdram_external_connection.local_refresh_ack
		output wire        local_wdata_req_from_the_ddr_sdram,   //                                         .local_wdata_req
		output wire        local_init_done_from_the_ddr_sdram,   //                                         .local_init_done
		output wire        reset_phy_clk_n_from_the_ddr_sdram,   //                                         .reset_phy_clk_n
		output wire        ddr_sdram_aux_half_rate_clk_out,      //                        ddr_sdram_auxhalf.clk
		output wire        ddr_sdram_aux_full_rate_clk_out,      //                        ddr_sdram_auxfull.clk
		input  wire        pll_areset_conduit_export,            //                       pll_areset_conduit.export
		output wire        pll_c2_out,                           //                               c2_out_clk.clk
		output wire        pll_c1_clk,                           //                                   pll_c1.clk
		output wire        pll_locked_conduit_export,            //                       pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export,         //                    pll_phasedone_conduit.export
		output wire        pll_c0_out,                           //                               c0_out_clk.clk
		output wire [1:0]  out_port_from_the_led_pio,            //              led_pio_external_connection.export
		input  wire [3:0]  in_port_to_the_button_pio,            //           button_pio_external_connection.export
		output wire        ddr_sdram_phy_clk_out,                //                           sysclk_out_clk.clk
		output wire [0:0]  read_n_to_the_ext_flash,              // flash_ssram_tristate_bridge_bridge_0_out.read_n_to_the_ext_flash
		output wire [0:0]  select_n_to_the_ext_flash,            //                                         .select_n_to_the_ext_flash
		output wire [23:0] flash_ssram_tristate_bridge_address,  //                                         .flash_ssram_tristate_bridge_address
		output wire [0:0]  bwe_n_to_the_ssram,                   //                                         .bwe_n_to_the_ssram
		output wire [0:0]  reset_n_to_the_ssram,                 //                                         .reset_n_to_the_ssram
		output wire [0:0]  chipenable1_n_to_the_ssram,           //                                         .chipenable1_n_to_the_ssram
		output wire [3:0]  bw_n_to_the_ssram,                    //                                         .bw_n_to_the_ssram
		output wire [0:0]  outputenable_n_to_the_ssram,          //                                         .outputenable_n_to_the_ssram
		inout  wire [31:0] flash_ssram_tristate_bridge_data,     //                                         .flash_ssram_tristate_bridge_data
		output wire [0:0]  adsc_n_to_the_ssram,                  //                                         .adsc_n_to_the_ssram
		output wire [0:0]  write_n_to_the_ext_flash,             //                                         .write_n_to_the_ext_flash
		inout  wire [0:0]  mem_clk_to_and_from_the_ddr_sdram,    //                         ddr_sdram_memory.mem_clk
		inout  wire [0:0]  mem_clk_n_to_and_from_the_ddr_sdram,  //                                         .mem_clk_n
		output wire [0:0]  mem_cs_n_from_the_ddr_sdram,          //                                         .mem_cs_n
		output wire [0:0]  mem_cke_from_the_ddr_sdram,           //                                         .mem_cke
		output wire [12:0] mem_addr_from_the_ddr_sdram,          //                                         .mem_addr
		output wire [1:0]  mem_ba_from_the_ddr_sdram,            //                                         .mem_ba
		output wire        mem_ras_n_from_the_ddr_sdram,         //                                         .mem_ras_n
		output wire        mem_cas_n_from_the_ddr_sdram,         //                                         .mem_cas_n
		output wire        mem_we_n_from_the_ddr_sdram,          //                                         .mem_we_n
		inout  wire [15:0] mem_dq_to_and_from_the_ddr_sdram,     //                                         .mem_dq
		inout  wire [1:0]  mem_dqs_to_and_from_the_ddr_sdram,    //                                         .mem_dqs
		output wire [1:0]  mem_dm_from_the_ddr_sdram,            //                                         .mem_dm
		input  wire        clk,                                  //                               clk_clk_in.clk
		input  wire        ddr_sdram_reset_n,                    //                 ddr_sdram_global_reset_n.reset_n
		output wire        pll_c3_out                            //                               c3_out_clk.clk
	);

	wire    [0:0] flash_ssram_pipeline_bridge_m0_burstcount;                                                              // flash_ssram_pipeline_bridge:m0_burstcount -> pipeline_bridge_before_tristate_bridge:s0_burstcount
	wire          flash_ssram_pipeline_bridge_m0_waitrequest;                                                             // pipeline_bridge_before_tristate_bridge:s0_waitrequest -> flash_ssram_pipeline_bridge:m0_waitrequest
	wire   [24:0] flash_ssram_pipeline_bridge_m0_address;                                                                 // flash_ssram_pipeline_bridge:m0_address -> pipeline_bridge_before_tristate_bridge:s0_address
	wire   [31:0] flash_ssram_pipeline_bridge_m0_writedata;                                                               // flash_ssram_pipeline_bridge:m0_writedata -> pipeline_bridge_before_tristate_bridge:s0_writedata
	wire          flash_ssram_pipeline_bridge_m0_write;                                                                   // flash_ssram_pipeline_bridge:m0_write -> pipeline_bridge_before_tristate_bridge:s0_write
	wire          flash_ssram_pipeline_bridge_m0_read;                                                                    // flash_ssram_pipeline_bridge:m0_read -> pipeline_bridge_before_tristate_bridge:s0_read
	wire   [31:0] flash_ssram_pipeline_bridge_m0_readdata;                                                                // pipeline_bridge_before_tristate_bridge:s0_readdata -> flash_ssram_pipeline_bridge:m0_readdata
	wire          flash_ssram_pipeline_bridge_m0_debugaccess;                                                             // flash_ssram_pipeline_bridge:m0_debugaccess -> pipeline_bridge_before_tristate_bridge:s0_debugaccess
	wire    [3:0] flash_ssram_pipeline_bridge_m0_byteenable;                                                              // flash_ssram_pipeline_bridge:m0_byteenable -> pipeline_bridge_before_tristate_bridge:s0_byteenable
	wire          flash_ssram_pipeline_bridge_m0_readdatavalid;                                                           // pipeline_bridge_before_tristate_bridge:s0_readdatavalid -> flash_ssram_pipeline_bridge:m0_readdatavalid
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out;                              // flash_ssram_tristate_bridge_pinSharer_0:select_n_to_the_ext_flash -> flash_ssram_tristate_bridge_bridge_0:tcs_select_n_to_the_ext_flash
	wire          flash_ssram_tristate_bridge_pinsharer_0_tcm_grant;                                                      // flash_ssram_tristate_bridge_bridge_0:grant -> flash_ssram_tristate_bridge_pinSharer_0:grant
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_outputenable_n_to_the_ssram_out;                            // flash_ssram_tristate_bridge_pinSharer_0:outputenable_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_outputenable_n_to_the_ssram
	wire   [31:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_in;                        // flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_data_in -> flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_data_in
	wire   [23:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_address_out;                    // flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_address -> flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_address
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out;                                // flash_ssram_tristate_bridge_pinSharer_0:read_n_to_the_ext_flash -> flash_ssram_tristate_bridge_bridge_0:tcs_read_n_to_the_ext_flash
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_adsc_n_to_the_ssram_out;                                    // flash_ssram_tristate_bridge_pinSharer_0:adsc_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_adsc_n_to_the_ssram
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out;                               // flash_ssram_tristate_bridge_pinSharer_0:write_n_to_the_ext_flash -> flash_ssram_tristate_bridge_bridge_0:tcs_write_n_to_the_ext_flash
	wire          flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_outen;                     // flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_data_outen -> flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_data_outen
	wire   [31:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_out;                       // flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_data -> flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_data
	wire          flash_ssram_tristate_bridge_pinsharer_0_tcm_request;                                                    // flash_ssram_tristate_bridge_pinSharer_0:request -> flash_ssram_tristate_bridge_bridge_0:request
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_bwe_n_to_the_ssram_out;                                     // flash_ssram_tristate_bridge_pinSharer_0:bwe_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_bwe_n_to_the_ssram
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_chipenable1_n_to_the_ssram_out;                             // flash_ssram_tristate_bridge_pinSharer_0:chipenable1_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_chipenable1_n_to_the_ssram
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_reset_n_to_the_ssram_out;                                   // flash_ssram_tristate_bridge_pinSharer_0:reset_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_reset_n_to_the_ssram
	wire    [3:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_bw_n_to_the_ssram_out;                                      // flash_ssram_tristate_bridge_pinSharer_0:bw_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_bw_n_to_the_ssram
	wire          ext_flash_tcm_chipselect_n_out;                                                                         // ext_flash:tcm_chipselect_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_chipselect_n_out
	wire          ext_flash_tcm_grant;                                                                                    // flash_ssram_tristate_bridge_pinSharer_0:tcs0_grant -> ext_flash:tcm_grant
	wire          ext_flash_tcm_data_outen;                                                                               // ext_flash:tcm_data_outen -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_data_outen
	wire          ext_flash_tcm_request;                                                                                  // ext_flash:tcm_request -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_request
	wire   [15:0] ext_flash_tcm_data_out;                                                                                 // ext_flash:tcm_data_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_data_out
	wire          ext_flash_tcm_write_n_out;                                                                              // ext_flash:tcm_write_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_write_n_out
	wire   [23:0] ext_flash_tcm_address_out;                                                                              // ext_flash:tcm_address_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_address_out
	wire   [15:0] ext_flash_tcm_data_in;                                                                                  // flash_ssram_tristate_bridge_pinSharer_0:tcs0_data_in -> ext_flash:tcm_data_in
	wire          ext_flash_tcm_read_n_out;                                                                               // ext_flash:tcm_read_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_read_n_out
	wire          ssram_tcm_chipselect_n_out;                                                                             // ssram:tcm_chipselect_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_chipselect_n_out
	wire          ssram_tcm_grant;                                                                                        // flash_ssram_tristate_bridge_pinSharer_0:tcs1_grant -> ssram:tcm_grant
	wire          ssram_tcm_data_outen;                                                                                   // ssram:tcm_data_outen -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_data_outen
	wire          ssram_tcm_reset_n_out;                                                                                  // ssram:tcm_reset_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_reset_n_out
	wire          ssram_tcm_outputenable_n_out;                                                                           // ssram:tcm_outputenable_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_outputenable_n_out
	wire          ssram_tcm_request;                                                                                      // ssram:tcm_request -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_request
	wire   [31:0] ssram_tcm_data_out;                                                                                     // ssram:tcm_data_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_data_out
	wire          ssram_tcm_write_n_out;                                                                                  // ssram:tcm_write_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_write_n_out
	wire   [19:0] ssram_tcm_address_out;                                                                                  // ssram:tcm_address_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_address_out
	wire   [31:0] ssram_tcm_data_in;                                                                                      // flash_ssram_tristate_bridge_pinSharer_0:tcs1_data_in -> ssram:tcm_data_in
	wire          ssram_tcm_begintransfer_n_out;                                                                          // ssram:tcm_begintransfer_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_begintransfer_n_out
	wire    [3:0] ssram_tcm_byteenable_n_out;                                                                             // ssram:tcm_byteenable_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_byteenable_n_out
	wire          cpu_data_master_waitrequest;                                                                            // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                              // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [27:0] cpu_data_master_address;                                                                                // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                  // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                   // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                               // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                            // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire          cpu_data_master_readdatavalid;                                                                          // cpu_data_master_translator:av_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                                                             // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          cpu_instruction_master_waitrequest;                                                                     // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [27:0] cpu_instruction_master_address;                                                                         // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                            // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                        // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                                   // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                         // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                           // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                        // cpu_jtag_debug_module_translator:av_chipselect -> cpu:jtag_debug_module_select
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                             // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                          // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                     // cpu_jtag_debug_module_translator:av_begintransfer -> cpu:jtag_debug_module_begintransfer
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                       // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                        // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                              // flash_ssram_pipeline_bridge:s0_waitrequest -> flash_ssram_pipeline_bridge_s0_translator:av_waitrequest
	wire    [0:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_burstcount;                               // flash_ssram_pipeline_bridge_s0_translator:av_burstcount -> flash_ssram_pipeline_bridge:s0_burstcount
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_writedata;                                // flash_ssram_pipeline_bridge_s0_translator:av_writedata -> flash_ssram_pipeline_bridge:s0_writedata
	wire   [24:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_address;                                  // flash_ssram_pipeline_bridge_s0_translator:av_address -> flash_ssram_pipeline_bridge:s0_address
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_write;                                    // flash_ssram_pipeline_bridge_s0_translator:av_write -> flash_ssram_pipeline_bridge:s0_write
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_read;                                     // flash_ssram_pipeline_bridge_s0_translator:av_read -> flash_ssram_pipeline_bridge:s0_read
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdata;                                 // flash_ssram_pipeline_bridge:s0_readdata -> flash_ssram_pipeline_bridge_s0_translator:av_readdata
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                              // flash_ssram_pipeline_bridge_s0_translator:av_debugaccess -> flash_ssram_pipeline_bridge:s0_debugaccess
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                            // flash_ssram_pipeline_bridge:s0_readdatavalid -> flash_ssram_pipeline_bridge_s0_translator:av_readdatavalid
	wire    [3:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_byteenable;                               // flash_ssram_pipeline_bridge_s0_translator:av_byteenable -> flash_ssram_pipeline_bridge:s0_byteenable
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                     // cpu_ddr_clock_bridge:s0_waitrequest -> cpu_ddr_clock_bridge_s0_translator:av_waitrequest
	wire    [0:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                      // cpu_ddr_clock_bridge_s0_translator:av_burstcount -> cpu_ddr_clock_bridge:s0_burstcount
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                       // cpu_ddr_clock_bridge_s0_translator:av_writedata -> cpu_ddr_clock_bridge:s0_writedata
	wire   [24:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                         // cpu_ddr_clock_bridge_s0_translator:av_address -> cpu_ddr_clock_bridge:s0_address
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                           // cpu_ddr_clock_bridge_s0_translator:av_write -> cpu_ddr_clock_bridge:s0_write
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                            // cpu_ddr_clock_bridge_s0_translator:av_read -> cpu_ddr_clock_bridge:s0_read
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                        // cpu_ddr_clock_bridge:s0_readdata -> cpu_ddr_clock_bridge_s0_translator:av_readdata
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                     // cpu_ddr_clock_bridge_s0_translator:av_debugaccess -> cpu_ddr_clock_bridge:s0_debugaccess
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                   // cpu_ddr_clock_bridge:s0_readdatavalid -> cpu_ddr_clock_bridge_s0_translator:av_readdatavalid
	wire    [3:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                      // cpu_ddr_clock_bridge_s0_translator:av_byteenable -> cpu_ddr_clock_bridge:s0_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                   // slow_peripheral_bridge:s0_waitrequest -> slow_peripheral_bridge_s0_translator:av_waitrequest
	wire    [0:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                    // slow_peripheral_bridge_s0_translator:av_burstcount -> slow_peripheral_bridge:s0_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata;                                     // slow_peripheral_bridge_s0_translator:av_writedata -> slow_peripheral_bridge:s0_writedata
	wire    [8:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address;                                       // slow_peripheral_bridge_s0_translator:av_address -> slow_peripheral_bridge:s0_address
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write;                                         // slow_peripheral_bridge_s0_translator:av_write -> slow_peripheral_bridge:s0_write
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read;                                          // slow_peripheral_bridge_s0_translator:av_read -> slow_peripheral_bridge:s0_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata;                                      // slow_peripheral_bridge:s0_readdata -> slow_peripheral_bridge_s0_translator:av_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                   // slow_peripheral_bridge_s0_translator:av_debugaccess -> slow_peripheral_bridge:s0_debugaccess
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                 // slow_peripheral_bridge:s0_readdatavalid -> slow_peripheral_bridge_s0_translator:av_readdatavalid
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                    // slow_peripheral_bridge_s0_translator:av_byteenable -> slow_peripheral_bridge:s0_byteenable
	wire    [0:0] cpu_ddr_clock_bridge_m0_burstcount;                                                                     // cpu_ddr_clock_bridge:m0_burstcount -> cpu_ddr_clock_bridge_m0_translator:av_burstcount
	wire          cpu_ddr_clock_bridge_m0_waitrequest;                                                                    // cpu_ddr_clock_bridge_m0_translator:av_waitrequest -> cpu_ddr_clock_bridge:m0_waitrequest
	wire   [24:0] cpu_ddr_clock_bridge_m0_address;                                                                        // cpu_ddr_clock_bridge:m0_address -> cpu_ddr_clock_bridge_m0_translator:av_address
	wire   [31:0] cpu_ddr_clock_bridge_m0_writedata;                                                                      // cpu_ddr_clock_bridge:m0_writedata -> cpu_ddr_clock_bridge_m0_translator:av_writedata
	wire          cpu_ddr_clock_bridge_m0_write;                                                                          // cpu_ddr_clock_bridge:m0_write -> cpu_ddr_clock_bridge_m0_translator:av_write
	wire          cpu_ddr_clock_bridge_m0_read;                                                                           // cpu_ddr_clock_bridge:m0_read -> cpu_ddr_clock_bridge_m0_translator:av_read
	wire   [31:0] cpu_ddr_clock_bridge_m0_readdata;                                                                       // cpu_ddr_clock_bridge_m0_translator:av_readdata -> cpu_ddr_clock_bridge:m0_readdata
	wire          cpu_ddr_clock_bridge_m0_debugaccess;                                                                    // cpu_ddr_clock_bridge:m0_debugaccess -> cpu_ddr_clock_bridge_m0_translator:av_debugaccess
	wire    [3:0] cpu_ddr_clock_bridge_m0_byteenable;                                                                     // cpu_ddr_clock_bridge:m0_byteenable -> cpu_ddr_clock_bridge_m0_translator:av_byteenable
	wire          cpu_ddr_clock_bridge_m0_readdatavalid;                                                                  // cpu_ddr_clock_bridge_m0_translator:av_readdatavalid -> cpu_ddr_clock_bridge:m0_readdatavalid
	wire          ddr_sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                // ddr_sdram:local_ready -> ddr_sdram_s1_translator:av_waitrequest
	wire    [0:0] ddr_sdram_s1_translator_avalon_anti_slave_0_burstcount;                                                 // ddr_sdram_s1_translator:av_burstcount -> ddr_sdram:local_size
	wire   [63:0] ddr_sdram_s1_translator_avalon_anti_slave_0_writedata;                                                  // ddr_sdram_s1_translator:av_writedata -> ddr_sdram:local_wdata
	wire   [21:0] ddr_sdram_s1_translator_avalon_anti_slave_0_address;                                                    // ddr_sdram_s1_translator:av_address -> ddr_sdram:local_address
	wire          ddr_sdram_s1_translator_avalon_anti_slave_0_write;                                                      // ddr_sdram_s1_translator:av_write -> ddr_sdram:local_write_req
	wire          ddr_sdram_s1_translator_avalon_anti_slave_0_beginbursttransfer;                                         // ddr_sdram_s1_translator:av_beginbursttransfer -> ddr_sdram:local_burstbegin
	wire          ddr_sdram_s1_translator_avalon_anti_slave_0_read;                                                       // ddr_sdram_s1_translator:av_read -> ddr_sdram:local_read_req
	wire   [63:0] ddr_sdram_s1_translator_avalon_anti_slave_0_readdata;                                                   // ddr_sdram:local_rdata -> ddr_sdram_s1_translator:av_readdata
	wire          ddr_sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                              // ddr_sdram:local_rdata_valid -> ddr_sdram_s1_translator:av_readdatavalid
	wire    [7:0] ddr_sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                 // ddr_sdram_s1_translator:av_byteenable -> ddr_sdram:local_be
	wire          ddr_sdram_reset_request_n_reset;                                                                        // ddr_sdram:reset_request_n -> [ddr_sdram_s1_translator:reset, ddr_sdram_s1_translator_avalon_universal_slave_0_agent:reset, ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_004:reset, rsp_xbar_demux_004:reset, rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1, width_adapter:reset, width_adapter_001:reset]
	wire    [0:0] slow_peripheral_bridge_m0_burstcount;                                                                   // slow_peripheral_bridge:m0_burstcount -> slow_peripheral_bridge_m0_translator:av_burstcount
	wire          slow_peripheral_bridge_m0_waitrequest;                                                                  // slow_peripheral_bridge_m0_translator:av_waitrequest -> slow_peripheral_bridge:m0_waitrequest
	wire    [8:0] slow_peripheral_bridge_m0_address;                                                                      // slow_peripheral_bridge:m0_address -> slow_peripheral_bridge_m0_translator:av_address
	wire   [31:0] slow_peripheral_bridge_m0_writedata;                                                                    // slow_peripheral_bridge:m0_writedata -> slow_peripheral_bridge_m0_translator:av_writedata
	wire          slow_peripheral_bridge_m0_write;                                                                        // slow_peripheral_bridge:m0_write -> slow_peripheral_bridge_m0_translator:av_write
	wire          slow_peripheral_bridge_m0_read;                                                                         // slow_peripheral_bridge:m0_read -> slow_peripheral_bridge_m0_translator:av_read
	wire   [31:0] slow_peripheral_bridge_m0_readdata;                                                                     // slow_peripheral_bridge_m0_translator:av_readdata -> slow_peripheral_bridge:m0_readdata
	wire          slow_peripheral_bridge_m0_debugaccess;                                                                  // slow_peripheral_bridge:m0_debugaccess -> slow_peripheral_bridge_m0_translator:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_byteenable;                                                                   // slow_peripheral_bridge:m0_byteenable -> slow_peripheral_bridge_m0_translator:av_byteenable
	wire          slow_peripheral_bridge_m0_readdatavalid;                                                                // slow_peripheral_bridge_m0_translator:av_readdatavalid -> slow_peripheral_bridge:m0_readdatavalid
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                                 // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire    [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                   // button_pio_s1_translator:av_address -> button_pio:address
	wire          button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire          button_pio_s1_translator_avalon_anti_slave_0_write;                                                     // button_pio_s1_translator:av_write -> button_pio:write_n
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire   [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_writedata;                                             // high_res_timer_s1_translator:av_writedata -> high_res_timer:writedata
	wire    [2:0] high_res_timer_s1_translator_avalon_anti_slave_0_address;                                               // high_res_timer_s1_translator:av_address -> high_res_timer:address
	wire          high_res_timer_s1_translator_avalon_anti_slave_0_chipselect;                                            // high_res_timer_s1_translator:av_chipselect -> high_res_timer:chipselect
	wire          high_res_timer_s1_translator_avalon_anti_slave_0_write;                                                 // high_res_timer_s1_translator:av_write -> high_res_timer:write_n
	wire   [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_readdata;                                              // high_res_timer:readdata -> high_res_timer_s1_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                 // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                   // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                     // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                  // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                       // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                        // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                    // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_writedata;                                                    // led_pio_s1_translator:av_writedata -> led_pio:writedata
	wire    [1:0] led_pio_s1_translator_avalon_anti_slave_0_address;                                                      // led_pio_s1_translator:av_address -> led_pio:address
	wire          led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led_pio_s1_translator:av_chipselect -> led_pio:chipselect
	wire          led_pio_s1_translator_avalon_anti_slave_0_write;                                                        // led_pio_s1_translator:av_write -> led_pio:write_n
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                     // led_pio:readdata -> led_pio_s1_translator:av_readdata
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_writedata;                             // performance_counter_control_slave_translator:av_writedata -> performance_counter:writedata
	wire    [2:0] performance_counter_control_slave_translator_avalon_anti_slave_0_address;                               // performance_counter_control_slave_translator:av_address -> performance_counter:address
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_write;                                 // performance_counter_control_slave_translator:av_write -> performance_counter:write
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_readdata;                              // performance_counter:readdata -> performance_counter_control_slave_translator:av_readdata
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer;                         // performance_counter_control_slave_translator:av_begintransfer -> performance_counter:begintransfer
	wire          remote_update_s1_translator_avalon_anti_slave_0_waitrequest;                                            // remote_update:waitrequest -> remote_update_s1_translator:av_waitrequest
	wire   [31:0] remote_update_s1_translator_avalon_anti_slave_0_writedata;                                              // remote_update_s1_translator:av_writedata -> remote_update:writedata
	wire    [5:0] remote_update_s1_translator_avalon_anti_slave_0_address;                                                // remote_update_s1_translator:av_address -> remote_update:address
	wire          remote_update_s1_translator_avalon_anti_slave_0_chipselect;                                             // remote_update_s1_translator:av_chipselect -> remote_update:chipselect
	wire          remote_update_s1_translator_avalon_anti_slave_0_write;                                                  // remote_update_s1_translator:av_write -> remote_update:write
	wire          remote_update_s1_translator_avalon_anti_slave_0_read;                                                   // remote_update_s1_translator:av_read -> remote_update:read
	wire   [31:0] remote_update_s1_translator_avalon_anti_slave_0_readdata;                                               // remote_update:readdata -> remote_update_s1_translator:av_readdata
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                              // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                                // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                             // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                                  // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                               // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                             // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                            // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_writedata;                                                 // pll_pll_slave_translator:av_writedata -> pll:writedata
	wire    [1:0] pll_pll_slave_translator_avalon_anti_slave_0_address;                                                   // pll_pll_slave_translator:av_address -> pll:address
	wire          pll_pll_slave_translator_avalon_anti_slave_0_write;                                                     // pll_pll_slave_translator:av_write -> pll:write
	wire          pll_pll_slave_translator_avalon_anti_slave_0_read;                                                      // pll_pll_slave_translator:av_read -> pll:read
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_readdata;                                                  // pll:readdata -> pll_pll_slave_translator:av_readdata
	wire    [0:0] pipeline_bridge_before_tristate_bridge_m0_burstcount;                                                   // pipeline_bridge_before_tristate_bridge:m0_burstcount -> pipeline_bridge_before_tristate_bridge_m0_translator:av_burstcount
	wire          pipeline_bridge_before_tristate_bridge_m0_waitrequest;                                                  // pipeline_bridge_before_tristate_bridge_m0_translator:av_waitrequest -> pipeline_bridge_before_tristate_bridge:m0_waitrequest
	wire   [24:0] pipeline_bridge_before_tristate_bridge_m0_address;                                                      // pipeline_bridge_before_tristate_bridge:m0_address -> pipeline_bridge_before_tristate_bridge_m0_translator:av_address
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_writedata;                                                    // pipeline_bridge_before_tristate_bridge:m0_writedata -> pipeline_bridge_before_tristate_bridge_m0_translator:av_writedata
	wire          pipeline_bridge_before_tristate_bridge_m0_write;                                                        // pipeline_bridge_before_tristate_bridge:m0_write -> pipeline_bridge_before_tristate_bridge_m0_translator:av_write
	wire          pipeline_bridge_before_tristate_bridge_m0_read;                                                         // pipeline_bridge_before_tristate_bridge:m0_read -> pipeline_bridge_before_tristate_bridge_m0_translator:av_read
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_readdata;                                                     // pipeline_bridge_before_tristate_bridge_m0_translator:av_readdata -> pipeline_bridge_before_tristate_bridge:m0_readdata
	wire          pipeline_bridge_before_tristate_bridge_m0_debugaccess;                                                  // pipeline_bridge_before_tristate_bridge:m0_debugaccess -> pipeline_bridge_before_tristate_bridge_m0_translator:av_debugaccess
	wire    [3:0] pipeline_bridge_before_tristate_bridge_m0_byteenable;                                                   // pipeline_bridge_before_tristate_bridge:m0_byteenable -> pipeline_bridge_before_tristate_bridge_m0_translator:av_byteenable
	wire          pipeline_bridge_before_tristate_bridge_m0_readdatavalid;                                                // pipeline_bridge_before_tristate_bridge_m0_translator:av_readdatavalid -> pipeline_bridge_before_tristate_bridge:m0_readdatavalid
	wire          ext_flash_uas_translator_avalon_anti_slave_0_waitrequest;                                               // ext_flash:uas_waitrequest -> ext_flash_uas_translator:av_waitrequest
	wire    [1:0] ext_flash_uas_translator_avalon_anti_slave_0_burstcount;                                                // ext_flash_uas_translator:av_burstcount -> ext_flash:uas_burstcount
	wire   [15:0] ext_flash_uas_translator_avalon_anti_slave_0_writedata;                                                 // ext_flash_uas_translator:av_writedata -> ext_flash:uas_writedata
	wire   [23:0] ext_flash_uas_translator_avalon_anti_slave_0_address;                                                   // ext_flash_uas_translator:av_address -> ext_flash:uas_address
	wire          ext_flash_uas_translator_avalon_anti_slave_0_lock;                                                      // ext_flash_uas_translator:av_lock -> ext_flash:uas_lock
	wire          ext_flash_uas_translator_avalon_anti_slave_0_write;                                                     // ext_flash_uas_translator:av_write -> ext_flash:uas_write
	wire          ext_flash_uas_translator_avalon_anti_slave_0_read;                                                      // ext_flash_uas_translator:av_read -> ext_flash:uas_read
	wire   [15:0] ext_flash_uas_translator_avalon_anti_slave_0_readdata;                                                  // ext_flash:uas_readdata -> ext_flash_uas_translator:av_readdata
	wire          ext_flash_uas_translator_avalon_anti_slave_0_debugaccess;                                               // ext_flash_uas_translator:av_debugaccess -> ext_flash:uas_debugaccess
	wire          ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid;                                             // ext_flash:uas_readdatavalid -> ext_flash_uas_translator:av_readdatavalid
	wire    [1:0] ext_flash_uas_translator_avalon_anti_slave_0_byteenable;                                                // ext_flash_uas_translator:av_byteenable -> ext_flash:uas_byteenable
	wire          ssram_uas_translator_avalon_anti_slave_0_waitrequest;                                                   // ssram:uas_waitrequest -> ssram_uas_translator:av_waitrequest
	wire    [2:0] ssram_uas_translator_avalon_anti_slave_0_burstcount;                                                    // ssram_uas_translator:av_burstcount -> ssram:uas_burstcount
	wire   [31:0] ssram_uas_translator_avalon_anti_slave_0_writedata;                                                     // ssram_uas_translator:av_writedata -> ssram:uas_writedata
	wire   [19:0] ssram_uas_translator_avalon_anti_slave_0_address;                                                       // ssram_uas_translator:av_address -> ssram:uas_address
	wire          ssram_uas_translator_avalon_anti_slave_0_lock;                                                          // ssram_uas_translator:av_lock -> ssram:uas_lock
	wire          ssram_uas_translator_avalon_anti_slave_0_write;                                                         // ssram_uas_translator:av_write -> ssram:uas_write
	wire          ssram_uas_translator_avalon_anti_slave_0_read;                                                          // ssram_uas_translator:av_read -> ssram:uas_read
	wire   [31:0] ssram_uas_translator_avalon_anti_slave_0_readdata;                                                      // ssram:uas_readdata -> ssram_uas_translator:av_readdata
	wire          ssram_uas_translator_avalon_anti_slave_0_debugaccess;                                                   // ssram_uas_translator:av_debugaccess -> ssram:uas_debugaccess
	wire          ssram_uas_translator_avalon_anti_slave_0_readdatavalid;                                                 // ssram:uas_readdatavalid -> ssram_uas_translator:av_readdatavalid
	wire    [3:0] ssram_uas_translator_avalon_anti_slave_0_byteenable;                                                    // ssram_uas_translator:av_byteenable -> ssram:uas_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                         // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_data_master_translator_avalon_universal_master_0_address;                                           // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                              // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                             // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                              // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                          // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                 // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                  // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [27:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                    // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                       // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                      // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                       // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                   // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                 // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [27:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                            // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // flash_ssram_pipeline_bridge_s0_translator:uav_waitrequest -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> flash_ssram_pipeline_bridge_s0_translator:uav_burstcount
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                  // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> flash_ssram_pipeline_bridge_s0_translator:uav_writedata
	wire   [27:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                    // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> flash_ssram_pipeline_bridge_s0_translator:uav_address
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                      // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> flash_ssram_pipeline_bridge_s0_translator:uav_write
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> flash_ssram_pipeline_bridge_s0_translator:uav_lock
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> flash_ssram_pipeline_bridge_s0_translator:uav_read
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                   // flash_ssram_pipeline_bridge_s0_translator:uav_readdata -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // flash_ssram_pipeline_bridge_s0_translator:uav_readdatavalid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> flash_ssram_pipeline_bridge_s0_translator:uav_debugaccess
	wire    [3:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> flash_ssram_pipeline_bridge_s0_translator:uav_byteenable
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;               // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;               // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // cpu_ddr_clock_bridge_s0_translator:uav_waitrequest -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_ddr_clock_bridge_s0_translator:uav_burstcount
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                         // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_ddr_clock_bridge_s0_translator:uav_writedata
	wire   [27:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                           // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_ddr_clock_bridge_s0_translator:uav_address
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                             // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_ddr_clock_bridge_s0_translator:uav_write
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                              // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_ddr_clock_bridge_s0_translator:uav_lock
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                              // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_ddr_clock_bridge_s0_translator:uav_read
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                          // cpu_ddr_clock_bridge_s0_translator:uav_readdata -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // cpu_ddr_clock_bridge_s0_translator:uav_readdatavalid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_ddr_clock_bridge_s0_translator:uav_debugaccess
	wire    [3:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_ddr_clock_bridge_s0_translator:uav_byteenable
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                       // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // slow_peripheral_bridge_s0_translator:uav_waitrequest -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> slow_peripheral_bridge_s0_translator:uav_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> slow_peripheral_bridge_s0_translator:uav_writedata
	wire   [27:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                         // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> slow_peripheral_bridge_s0_translator:uav_address
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> slow_peripheral_bridge_s0_translator:uav_write
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> slow_peripheral_bridge_s0_translator:uav_lock
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> slow_peripheral_bridge_s0_translator:uav_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // slow_peripheral_bridge_s0_translator:uav_readdata -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // slow_peripheral_bridge_s0_translator:uav_readdatavalid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> slow_peripheral_bridge_s0_translator:uav_debugaccess
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> slow_peripheral_bridge_s0_translator:uav_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [99:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [99:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                               // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_ddr_clock_bridge_m0_translator:uav_waitrequest
	wire    [2:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                                // cpu_ddr_clock_bridge_m0_translator:uav_burstcount -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                 // cpu_ddr_clock_bridge_m0_translator:uav_writedata -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address;                                   // cpu_ddr_clock_bridge_m0_translator:uav_address -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                      // cpu_ddr_clock_bridge_m0_translator:uav_lock -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write;                                     // cpu_ddr_clock_bridge_m0_translator:uav_write -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read;                                      // cpu_ddr_clock_bridge_m0_translator:uav_read -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                  // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_ddr_clock_bridge_m0_translator:uav_readdata
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                               // cpu_ddr_clock_bridge_m0_translator:uav_debugaccess -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                                // cpu_ddr_clock_bridge_m0_translator:uav_byteenable -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                             // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_ddr_clock_bridge_m0_translator:uav_readdatavalid
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // ddr_sdram_s1_translator:uav_waitrequest -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [3:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr_sdram_s1_translator:uav_burstcount
	wire   [63:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr_sdram_s1_translator:uav_writedata
	wire   [24:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr_sdram_s1_translator:uav_address
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr_sdram_s1_translator:uav_write
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr_sdram_s1_translator:uav_lock
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr_sdram_s1_translator:uav_read
	wire   [63:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // ddr_sdram_s1_translator:uav_readdata -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // ddr_sdram_s1_translator:uav_readdatavalid -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr_sdram_s1_translator:uav_debugaccess
	wire    [7:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr_sdram_s1_translator:uav_byteenable
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [132:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [132:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [63:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest;                             // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> slow_peripheral_bridge_m0_translator:uav_waitrequest
	wire    [2:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount;                              // slow_peripheral_bridge_m0_translator:uav_burstcount -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata;                               // slow_peripheral_bridge_m0_translator:uav_writedata -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [8:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address;                                 // slow_peripheral_bridge_m0_translator:uav_address -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock;                                    // slow_peripheral_bridge_m0_translator:uav_lock -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write;                                   // slow_peripheral_bridge_m0_translator:uav_write -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read;                                    // slow_peripheral_bridge_m0_translator:uav_read -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata;                                // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> slow_peripheral_bridge_m0_translator:uav_readdata
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess;                             // slow_peripheral_bridge_m0_translator:uav_debugaccess -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable;                              // slow_peripheral_bridge_m0_translator:uav_byteenable -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                           // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> slow_peripheral_bridge_m0_translator:uav_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire    [8:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire    [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // high_res_timer_s1_translator:uav_waitrequest -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_res_timer_s1_translator:uav_burstcount
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_res_timer_s1_translator:uav_writedata
	wire    [8:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_res_timer_s1_translator:uav_address
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_res_timer_s1_translator:uav_write
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_res_timer_s1_translator:uav_lock
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_res_timer_s1_translator:uav_read
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // high_res_timer_s1_translator:uav_readdata -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // high_res_timer_s1_translator:uav_readdatavalid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_res_timer_s1_translator:uav_debugaccess
	wire    [3:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_res_timer_s1_translator:uav_byteenable
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire    [8:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led_pio_s1_translator:uav_waitrequest -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_pio_s1_translator:uav_burstcount
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_pio_s1_translator:uav_writedata
	wire    [8:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_pio_s1_translator:uav_address
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_pio_s1_translator:uav_write
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_pio_s1_translator:uav_lock
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_pio_s1_translator:uav_read
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led_pio_s1_translator:uav_readdata -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led_pio_s1_translator:uav_readdatavalid -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_pio_s1_translator:uav_debugaccess
	wire    [3:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_pio_s1_translator:uav_byteenable
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // performance_counter_control_slave_translator:uav_waitrequest -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_control_slave_translator:uav_burstcount
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_control_slave_translator:uav_writedata
	wire    [8:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_control_slave_translator:uav_address
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_control_slave_translator:uav_write
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_control_slave_translator:uav_lock
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_control_slave_translator:uav_read
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // performance_counter_control_slave_translator:uav_readdata -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // performance_counter_control_slave_translator:uav_readdatavalid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_control_slave_translator:uav_debugaccess
	wire    [3:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_control_slave_translator:uav_byteenable
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // remote_update_s1_translator:uav_waitrequest -> remote_update_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] remote_update_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> remote_update_s1_translator:uav_burstcount
	wire   [31:0] remote_update_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> remote_update_s1_translator:uav_writedata
	wire    [8:0] remote_update_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_address -> remote_update_s1_translator:uav_address
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_write -> remote_update_s1_translator:uav_write
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_lock -> remote_update_s1_translator:uav_lock
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_read -> remote_update_s1_translator:uav_read
	wire   [31:0] remote_update_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // remote_update_s1_translator:uav_readdata -> remote_update_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // remote_update_s1_translator:uav_readdatavalid -> remote_update_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> remote_update_s1_translator:uav_debugaccess
	wire    [3:0] remote_update_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // remote_update_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> remote_update_s1_translator:uav_byteenable
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // remote_update_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // remote_update_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // remote_update_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // remote_update_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> remote_update_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> remote_update_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> remote_update_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> remote_update_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> remote_update_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // remote_update_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // remote_update_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // remote_update_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> remote_update_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> remote_update_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> remote_update_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // remote_update_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire    [8:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [8:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // pll_pll_slave_translator:uav_waitrequest -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pll_pll_slave_translator:uav_burstcount
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pll_pll_slave_translator:uav_writedata
	wire    [8:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                     // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> pll_pll_slave_translator:uav_address
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> pll_pll_slave_translator:uav_write
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pll_pll_slave_translator:uav_lock
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> pll_pll_slave_translator:uav_read
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // pll_pll_slave_translator:uav_readdata -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // pll_pll_slave_translator:uav_readdatavalid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pll_pll_slave_translator:uav_debugaccess
	wire    [3:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pll_pll_slave_translator:uav_byteenable
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_waitrequest;             // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> pipeline_bridge_before_tristate_bridge_m0_translator:uav_waitrequest
	wire    [2:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_burstcount;              // pipeline_bridge_before_tristate_bridge_m0_translator:uav_burstcount -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_writedata;               // pipeline_bridge_before_tristate_bridge_m0_translator:uav_writedata -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_address;                 // pipeline_bridge_before_tristate_bridge_m0_translator:uav_address -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_lock;                    // pipeline_bridge_before_tristate_bridge_m0_translator:uav_lock -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_write;                   // pipeline_bridge_before_tristate_bridge_m0_translator:uav_write -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_read;                    // pipeline_bridge_before_tristate_bridge_m0_translator:uav_read -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdata;                // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> pipeline_bridge_before_tristate_bridge_m0_translator:uav_readdata
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_debugaccess;             // pipeline_bridge_before_tristate_bridge_m0_translator:uav_debugaccess -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_byteenable;              // pipeline_bridge_before_tristate_bridge_m0_translator:uav_byteenable -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdatavalid;           // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> pipeline_bridge_before_tristate_bridge_m0_translator:uav_readdatavalid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // ext_flash_uas_translator:uav_waitrequest -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> ext_flash_uas_translator:uav_burstcount
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> ext_flash_uas_translator:uav_writedata
	wire   [24:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address;                                     // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_address -> ext_flash_uas_translator:uav_address
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write;                                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_write -> ext_flash_uas_translator:uav_write
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_lock -> ext_flash_uas_translator:uav_lock
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_read -> ext_flash_uas_translator:uav_read
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // ext_flash_uas_translator:uav_readdata -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // ext_flash_uas_translator:uav_readdatavalid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ext_flash_uas_translator:uav_debugaccess
	wire    [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> ext_flash_uas_translator:uav_byteenable
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [76:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [76:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // ssram_uas_translator:uav_waitrequest -> ssram_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // ssram_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> ssram_uas_translator:uav_burstcount
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // ssram_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> ssram_uas_translator:uav_writedata
	wire   [24:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_address;                                         // ssram_uas_translator_avalon_universal_slave_0_agent:m0_address -> ssram_uas_translator:uav_address
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_write;                                           // ssram_uas_translator_avalon_universal_slave_0_agent:m0_write -> ssram_uas_translator:uav_write
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                            // ssram_uas_translator_avalon_universal_slave_0_agent:m0_lock -> ssram_uas_translator:uav_lock
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_read;                                            // ssram_uas_translator_avalon_universal_slave_0_agent:m0_read -> ssram_uas_translator:uav_read
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // ssram_uas_translator:uav_readdata -> ssram_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // ssram_uas_translator:uav_readdatavalid -> ssram_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // ssram_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ssram_uas_translator:uav_debugaccess
	wire    [3:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // ssram_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> ssram_uas_translator:uav_byteenable
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [94:0] ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [94:0] ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [98:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [98:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_001:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire   [98:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                      // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [98:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_001:sink_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                             // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [98:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                              // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_002:sink_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [98:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_003:sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                            // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [95:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                             // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_002:sink_ready -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [131:0] ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_004:sink_ready -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                    // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                          // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                  // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [83:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                           // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                          // addr_router_003:sink_ready -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [83:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_005:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [83:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_006:sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_007:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [83:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_008:sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [83:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_009:sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // remote_update_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // remote_update_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // remote_update_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [83:0] remote_update_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // remote_update_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          remote_update_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_010:sink_ready -> remote_update_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [83:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_011:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [83:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_012:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [83:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_013:sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;    // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;          // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;  // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [93:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;           // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;          // addr_router_004:sink_ready -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [75:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_014:sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // ssram_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                           // ssram_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // ssram_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [93:0] ssram_uas_translator_avalon_universal_slave_0_agent_rp_data;                                            // ssram_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_015:sink_ready -> ssram_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire   [98:0] addr_router_src_data;                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire    [3:0] addr_router_src_channel;                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                            // limiter:rsp_src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                  // limiter:rsp_src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                          // limiter:rsp_src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [98:0] limiter_rsp_src_data;                                                                                   // limiter:rsp_src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] limiter_rsp_src_channel;                                                                                // limiter:rsp_src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                  // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                        // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                              // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                      // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [98:0] addr_router_001_src_data;                                                                               // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire    [3:0] addr_router_001_src_channel;                                                                            // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                              // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                        // limiter_001:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                              // limiter_001:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                      // limiter_001:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [98:0] limiter_001_rsp_src_data;                                                                               // limiter_001:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] limiter_001_rsp_src_channel;                                                                            // limiter_001:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_003_src_endofpacket;                                                                        // addr_router_003:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                              // addr_router_003:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                      // addr_router_003:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [83:0] addr_router_003_src_data;                                                                               // addr_router_003:src_data -> limiter_002:cmd_sink_data
	wire    [8:0] addr_router_003_src_channel;                                                                            // addr_router_003:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                              // limiter_002:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                        // limiter_002:rsp_src_endofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                              // limiter_002:rsp_src_valid -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                      // limiter_002:rsp_src_startofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [83:0] limiter_002_rsp_src_data;                                                                               // limiter_002:rsp_src_data -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [8:0] limiter_002_rsp_src_channel;                                                                            // limiter_002:rsp_src_channel -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                              // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          addr_router_004_src_endofpacket;                                                                        // addr_router_004:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire          addr_router_004_src_valid;                                                                              // addr_router_004:src_valid -> limiter_003:cmd_sink_valid
	wire          addr_router_004_src_startofpacket;                                                                      // addr_router_004:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire   [93:0] addr_router_004_src_data;                                                                               // addr_router_004:src_data -> limiter_003:cmd_sink_data
	wire    [1:0] addr_router_004_src_channel;                                                                            // addr_router_004:src_channel -> limiter_003:cmd_sink_channel
	wire          addr_router_004_src_ready;                                                                              // limiter_003:cmd_sink_ready -> addr_router_004:src_ready
	wire          limiter_003_rsp_src_endofpacket;                                                                        // limiter_003:rsp_src_endofpacket -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_003_rsp_src_valid;                                                                              // limiter_003:rsp_src_valid -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_003_rsp_src_startofpacket;                                                                      // limiter_003:rsp_src_startofpacket -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [93:0] limiter_003_rsp_src_data;                                                                               // limiter_003:rsp_src_data -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] limiter_003_rsp_src_channel;                                                                            // limiter_003:rsp_src_channel -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_003_rsp_src_ready;                                                                              // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                      // burst_adapter:source0_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                            // burst_adapter:source0_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                    // burst_adapter:source0_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [75:0] burst_adapter_source0_data;                                                                             // burst_adapter:source0_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                                          // burst_adapter:source0_channel -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                         // rst_controller:reset_out -> ddr_sdram:soft_reset_n
	wire          cpu_jtag_debug_module_reset_reset;                                                                      // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2, rst_controller_004:reset_in2]
	wire          rst_controller_001_reset_out_reset;                                                                     // rst_controller_001:reset_out -> [addr_router_003:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_003:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, high_res_timer:reset_n, high_res_timer_s1_translator:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_011:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_pio:reset_n, led_pio_s1_translator:reset, led_pio_s1_translator_avalon_universal_slave_0_agent:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, performance_counter:reset_n, performance_counter_control_slave_translator:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_011:reset, rsp_xbar_mux_003:reset, slow_peripheral_bridge:m0_reset, slow_peripheral_bridge_m0_translator:reset, slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_002_reset_out_reset;                                                                     // rst_controller_002:reset_out -> [crosser:out_reset, crosser_003:in_reset, id_router_010:reset, remote_update:reset, remote_update_s1_translator:reset, remote_update_s1_translator_avalon_universal_slave_0_agent:reset, remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_010:reset]
	wire          rst_controller_003_reset_out_reset;                                                                     // rst_controller_003:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_004:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_ddr_clock_bridge:s0_reset, cpu_ddr_clock_bridge_s0_translator:reset, cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser_001:out_reset, crosser_004:in_reset, ext_flash:reset_reset, ext_flash_uas_translator:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_ssram_pipeline_bridge:reset, flash_ssram_pipeline_bridge_s0_translator:reset, flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:reset, flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_ssram_tristate_bridge_bridge_0:reset, flash_ssram_tristate_bridge_pinSharer_0:reset_reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_012:reset, id_router_014:reset, id_router_015:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, limiter:reset, limiter_001:reset, limiter_003:reset, pipeline_bridge_before_tristate_bridge:reset, pipeline_bridge_before_tristate_bridge_m0_translator:reset, pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_004:reset, slow_peripheral_bridge:s0_reset, slow_peripheral_bridge_s0_translator:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ssram:reset_reset, ssram_uas_translator:reset, ssram_uas_translator_avalon_universal_slave_0_agent:reset, ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_004_reset_out_reset;                                                                     // rst_controller_004:reset_out -> [addr_router_002:reset, cmd_xbar_demux_002:reset, cpu_ddr_clock_bridge:m0_reset, cpu_ddr_clock_bridge_m0_translator:reset, cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset]
	wire          rst_controller_005_reset_out_reset;                                                                     // rst_controller_005:reset_out -> [crosser_002:out_reset, crosser_005:in_reset, id_router_013:reset, pll:reset, pll_pll_slave_translator:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_013:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                        // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                              // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                      // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire   [98:0] cmd_xbar_demux_src0_data;                                                                               // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [3:0] cmd_xbar_demux_src0_channel;                                                                            // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                              // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                        // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                              // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                      // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [98:0] cmd_xbar_demux_src1_data;                                                                               // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [3:0] cmd_xbar_demux_src1_channel;                                                                            // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                              // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                        // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                              // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                      // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [98:0] cmd_xbar_demux_src2_data;                                                                               // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire    [3:0] cmd_xbar_demux_src2_channel;                                                                            // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                              // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                        // cmd_xbar_demux:src3_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                              // cmd_xbar_demux:src3_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                      // cmd_xbar_demux:src3_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] cmd_xbar_demux_src3_data;                                                                               // cmd_xbar_demux:src3_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_demux_src3_channel;                                                                            // cmd_xbar_demux:src3_channel -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                    // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                          // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                  // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire   [98:0] cmd_xbar_demux_001_src0_data;                                                                           // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [3:0] cmd_xbar_demux_001_src0_channel;                                                                        // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                          // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                    // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                          // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                  // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [98:0] cmd_xbar_demux_001_src1_data;                                                                           // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [3:0] cmd_xbar_demux_001_src1_channel;                                                                        // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                          // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                    // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                          // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                  // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [98:0] cmd_xbar_demux_001_src2_data;                                                                           // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire    [3:0] cmd_xbar_demux_001_src2_channel;                                                                        // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                          // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [98:0] rsp_xbar_demux_src0_data;                                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [3:0] rsp_xbar_demux_src0_channel;                                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                        // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                              // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                      // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire   [98:0] rsp_xbar_demux_src1_data;                                                                               // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [3:0] rsp_xbar_demux_src1_channel;                                                                            // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                              // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [98:0] rsp_xbar_demux_001_src0_data;                                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [3:0] rsp_xbar_demux_001_src0_channel;                                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                    // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                          // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                  // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire   [98:0] rsp_xbar_demux_001_src1_data;                                                                           // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [3:0] rsp_xbar_demux_001_src1_channel;                                                                        // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                          // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire   [98:0] rsp_xbar_demux_002_src0_data;                                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [3:0] rsp_xbar_demux_002_src0_channel;                                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                    // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                          // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                  // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire   [98:0] rsp_xbar_demux_002_src1_data;                                                                           // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire    [3:0] rsp_xbar_demux_002_src1_channel;                                                                        // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                          // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire   [98:0] rsp_xbar_demux_003_src0_data;                                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [3:0] rsp_xbar_demux_003_src0_channel;                                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                          // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [98:0] limiter_cmd_src_data;                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [3:0] limiter_cmd_src_channel;                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire   [98:0] rsp_xbar_mux_src_data;                                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [3:0] rsp_xbar_mux_src_channel;                                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                        // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                      // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [98:0] limiter_001_cmd_src_data;                                                                               // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire    [3:0] limiter_001_cmd_src_channel;                                                                            // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                              // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                       // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                             // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                     // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [98:0] rsp_xbar_mux_001_src_data;                                                                              // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire    [3:0] rsp_xbar_mux_001_src_channel;                                                                           // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                             // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                           // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                 // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                         // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] cmd_xbar_mux_src_data;                                                                                  // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_src_channel;                                                                               // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [98:0] id_router_src_data;                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [3:0] id_router_src_channel;                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                       // cmd_xbar_mux_001:src_endofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                             // cmd_xbar_mux_001:src_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                     // cmd_xbar_mux_001:src_startofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] cmd_xbar_mux_001_src_data;                                                                              // cmd_xbar_mux_001:src_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_001_src_channel;                                                                           // cmd_xbar_mux_001:src_channel -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                             // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [98:0] id_router_001_src_data;                                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [3:0] id_router_001_src_channel;                                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                       // cmd_xbar_mux_002:src_endofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                             // cmd_xbar_mux_002:src_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                     // cmd_xbar_mux_002:src_startofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [98:0] cmd_xbar_mux_002_src_data;                                                                              // cmd_xbar_mux_002:src_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_002_src_channel;                                                                           // cmd_xbar_mux_002:src_channel -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                             // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [98:0] id_router_002_src_data;                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [3:0] id_router_002_src_channel;                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_src3_ready;                                                                              // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire          id_router_003_src_endofpacket;                                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [98:0] id_router_003_src_data;                                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [3:0] id_router_003_src_channel;                                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                    // cmd_xbar_demux_002:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                          // cmd_xbar_demux_002:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                  // cmd_xbar_demux_002:src0_startofpacket -> width_adapter:in_startofpacket
	wire   [95:0] cmd_xbar_demux_002_src0_data;                                                                           // cmd_xbar_demux_002:src0_data -> width_adapter:in_data
	wire    [0:0] cmd_xbar_demux_002_src0_channel;                                                                        // cmd_xbar_demux_002:src0_channel -> width_adapter:in_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                    // rsp_xbar_demux_004:src0_endofpacket -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                          // rsp_xbar_demux_004:src0_valid -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                  // rsp_xbar_demux_004:src0_startofpacket -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [95:0] rsp_xbar_demux_004_src0_data;                                                                           // rsp_xbar_demux_004:src0_data -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_004_src0_channel;                                                                        // rsp_xbar_demux_004:src0_channel -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_002_src_endofpacket;                                                                        // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                              // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                      // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [95:0] addr_router_002_src_data;                                                                               // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [0:0] addr_router_002_src_channel;                                                                            // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                              // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_004_src0_ready;                                                                          // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                    // cmd_xbar_demux_003:src0_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                          // cmd_xbar_demux_003:src0_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                  // cmd_xbar_demux_003:src0_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src0_data;                                                                           // cmd_xbar_demux_003:src0_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_003_src0_channel;                                                                        // cmd_xbar_demux_003:src0_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                    // cmd_xbar_demux_003:src1_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                          // cmd_xbar_demux_003:src1_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                                  // cmd_xbar_demux_003:src1_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src1_data;                                                                           // cmd_xbar_demux_003:src1_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_003_src1_channel;                                                                        // cmd_xbar_demux_003:src1_channel -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src2_endofpacket;                                                                    // cmd_xbar_demux_003:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src2_valid;                                                                          // cmd_xbar_demux_003:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src2_startofpacket;                                                                  // cmd_xbar_demux_003:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src2_data;                                                                           // cmd_xbar_demux_003:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_003_src2_channel;                                                                        // cmd_xbar_demux_003:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src3_endofpacket;                                                                    // cmd_xbar_demux_003:src3_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src3_valid;                                                                          // cmd_xbar_demux_003:src3_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src3_startofpacket;                                                                  // cmd_xbar_demux_003:src3_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src3_data;                                                                           // cmd_xbar_demux_003:src3_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_003_src3_channel;                                                                        // cmd_xbar_demux_003:src3_channel -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src4_endofpacket;                                                                    // cmd_xbar_demux_003:src4_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src4_valid;                                                                          // cmd_xbar_demux_003:src4_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src4_startofpacket;                                                                  // cmd_xbar_demux_003:src4_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src4_data;                                                                           // cmd_xbar_demux_003:src4_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_003_src4_channel;                                                                        // cmd_xbar_demux_003:src4_channel -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src6_endofpacket;                                                                    // cmd_xbar_demux_003:src6_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src6_valid;                                                                          // cmd_xbar_demux_003:src6_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src6_startofpacket;                                                                  // cmd_xbar_demux_003:src6_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src6_data;                                                                           // cmd_xbar_demux_003:src6_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] cmd_xbar_demux_003_src6_channel;                                                                        // cmd_xbar_demux_003:src6_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                    // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                          // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                  // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire   [83:0] rsp_xbar_demux_005_src0_data;                                                                           // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_003:sink0_data
	wire    [8:0] rsp_xbar_demux_005_src0_channel;                                                                        // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                          // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire   [83:0] rsp_xbar_demux_006_src0_data;                                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_003:sink1_data
	wire    [8:0] rsp_xbar_demux_006_src0_channel;                                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                          // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_003:sink2_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire   [83:0] rsp_xbar_demux_007_src0_data;                                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_003:sink2_data
	wire    [8:0] rsp_xbar_demux_007_src0_channel;                                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_003:sink2_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                          // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                    // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_003:sink3_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                          // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_003:sink3_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                  // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_003:sink3_startofpacket
	wire   [83:0] rsp_xbar_demux_008_src0_data;                                                                           // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_003:sink3_data
	wire    [8:0] rsp_xbar_demux_008_src0_channel;                                                                        // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_003:sink3_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                          // rsp_xbar_mux_003:sink3_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                    // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_003:sink4_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                          // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_003:sink4_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                  // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_003:sink4_startofpacket
	wire   [83:0] rsp_xbar_demux_009_src0_data;                                                                           // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_003:sink4_data
	wire    [8:0] rsp_xbar_demux_009_src0_channel;                                                                        // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_003:sink4_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                          // rsp_xbar_mux_003:sink4_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                    // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_003:sink6_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                          // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_003:sink6_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                  // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_003:sink6_startofpacket
	wire   [83:0] rsp_xbar_demux_011_src0_data;                                                                           // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_003:sink6_data
	wire    [8:0] rsp_xbar_demux_011_src0_channel;                                                                        // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_003:sink6_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                          // rsp_xbar_mux_003:sink6_ready -> rsp_xbar_demux_011:src0_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                        // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                      // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [83:0] limiter_002_cmd_src_data;                                                                               // limiter_002:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire    [8:0] limiter_002_cmd_src_channel;                                                                            // limiter_002:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                              // cmd_xbar_demux_003:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                       // rsp_xbar_mux_003:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                             // rsp_xbar_mux_003:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                     // rsp_xbar_mux_003:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [83:0] rsp_xbar_mux_003_src_data;                                                                              // rsp_xbar_mux_003:src_data -> limiter_002:rsp_sink_data
	wire    [8:0] rsp_xbar_mux_003_src_channel;                                                                           // rsp_xbar_mux_003:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                             // limiter_002:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          cmd_xbar_demux_003_src0_ready;                                                                          // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src0_ready
	wire          id_router_005_src_endofpacket;                                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [83:0] id_router_005_src_data;                                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [8:0] id_router_005_src_channel;                                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_003_src1_ready;                                                                          // high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src1_ready
	wire          id_router_006_src_endofpacket;                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [83:0] id_router_006_src_data;                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [8:0] id_router_006_src_channel;                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_003_src2_ready;                                                                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src2_ready
	wire          id_router_007_src_endofpacket;                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [83:0] id_router_007_src_data;                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [8:0] id_router_007_src_channel;                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_003_src3_ready;                                                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src3_ready
	wire          id_router_008_src_endofpacket;                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [83:0] id_router_008_src_data;                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [8:0] id_router_008_src_channel;                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_003_src4_ready;                                                                          // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src4_ready
	wire          id_router_009_src_endofpacket;                                                                          // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                        // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [83:0] id_router_009_src_data;                                                                                 // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire    [8:0] id_router_009_src_channel;                                                                              // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          crosser_out_ready;                                                                                      // remote_update_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_010_src_endofpacket;                                                                          // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                        // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [83:0] id_router_010_src_data;                                                                                 // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire    [8:0] id_router_010_src_channel;                                                                              // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_003_src6_ready;                                                                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src6_ready
	wire          id_router_011_src_endofpacket;                                                                          // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                        // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [83:0] id_router_011_src_data;                                                                                 // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire    [8:0] id_router_011_src_channel;                                                                              // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          crosser_001_out_ready;                                                                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire          id_router_012_src_endofpacket;                                                                          // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                        // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [83:0] id_router_012_src_data;                                                                                 // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire    [8:0] id_router_012_src_channel;                                                                              // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          crosser_002_out_ready;                                                                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire          id_router_013_src_endofpacket;                                                                          // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                        // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [83:0] id_router_013_src_data;                                                                                 // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire    [8:0] id_router_013_src_channel;                                                                              // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                    // cmd_xbar_demux_004:src0_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                          // cmd_xbar_demux_004:src0_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                  // cmd_xbar_demux_004:src0_startofpacket -> width_adapter_002:in_startofpacket
	wire   [93:0] cmd_xbar_demux_004_src0_data;                                                                           // cmd_xbar_demux_004:src0_data -> width_adapter_002:in_data
	wire    [1:0] cmd_xbar_demux_004_src0_channel;                                                                        // cmd_xbar_demux_004:src0_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                                    // cmd_xbar_demux_004:src1_endofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                          // cmd_xbar_demux_004:src1_valid -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                                  // cmd_xbar_demux_004:src1_startofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [93:0] cmd_xbar_demux_004_src1_data;                                                                           // cmd_xbar_demux_004:src1_data -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] cmd_xbar_demux_004_src1_channel;                                                                        // cmd_xbar_demux_004:src1_channel -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                    // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                          // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_004:sink0_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                  // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire   [93:0] rsp_xbar_demux_014_src0_data;                                                                           // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_004:sink0_data
	wire    [1:0] rsp_xbar_demux_014_src0_channel;                                                                        // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_004:sink0_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                          // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                    // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                          // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_004:sink1_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                  // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire   [93:0] rsp_xbar_demux_015_src0_data;                                                                           // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_004:sink1_data
	wire    [1:0] rsp_xbar_demux_015_src0_channel;                                                                        // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_004:sink1_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                          // rsp_xbar_mux_004:sink1_ready -> rsp_xbar_demux_015:src0_ready
	wire          limiter_003_cmd_src_endofpacket;                                                                        // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          limiter_003_cmd_src_startofpacket;                                                                      // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [93:0] limiter_003_cmd_src_data;                                                                               // limiter_003:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire    [1:0] limiter_003_cmd_src_channel;                                                                            // limiter_003:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire          limiter_003_cmd_src_ready;                                                                              // cmd_xbar_demux_004:sink_ready -> limiter_003:cmd_src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                       // rsp_xbar_mux_004:src_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                             // rsp_xbar_mux_004:src_valid -> limiter_003:rsp_sink_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                                     // rsp_xbar_mux_004:src_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire   [93:0] rsp_xbar_mux_004_src_data;                                                                              // rsp_xbar_mux_004:src_data -> limiter_003:rsp_sink_data
	wire    [1:0] rsp_xbar_mux_004_src_channel;                                                                           // rsp_xbar_mux_004:src_channel -> limiter_003:rsp_sink_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                             // limiter_003:rsp_sink_ready -> rsp_xbar_mux_004:src_ready
	wire          cmd_xbar_demux_004_src1_ready;                                                                          // ssram_uas_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src1_ready
	wire          id_router_015_src_endofpacket;                                                                          // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                        // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [93:0] id_router_015_src_data;                                                                                 // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire    [1:0] id_router_015_src_channel;                                                                              // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_002_src0_ready;                                                                          // width_adapter:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          width_adapter_src_endofpacket;                                                                          // width_adapter:out_endofpacket -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          width_adapter_src_valid;                                                                                // width_adapter:out_valid -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          width_adapter_src_startofpacket;                                                                        // width_adapter:out_startofpacket -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [131:0] width_adapter_src_data;                                                                                 // width_adapter:out_data -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          width_adapter_src_ready;                                                                                // ddr_sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter:out_ready
	wire          width_adapter_src_channel;                                                                              // width_adapter:out_channel -> ddr_sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          id_router_004_src_endofpacket;                                                                          // id_router_004:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_004_src_valid;                                                                                // id_router_004:src_valid -> width_adapter_001:in_valid
	wire          id_router_004_src_startofpacket;                                                                        // id_router_004:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [131:0] id_router_004_src_data;                                                                                 // id_router_004:src_data -> width_adapter_001:in_data
	wire    [0:0] id_router_004_src_channel;                                                                              // id_router_004:src_channel -> width_adapter_001:in_channel
	wire          id_router_004_src_ready;                                                                                // width_adapter_001:in_ready -> id_router_004:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                      // width_adapter_001:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                            // width_adapter_001:out_valid -> rsp_xbar_demux_004:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                    // width_adapter_001:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [95:0] width_adapter_001_src_data;                                                                             // width_adapter_001:out_data -> rsp_xbar_demux_004:sink_data
	wire          width_adapter_001_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> width_adapter_001:out_ready
	wire          width_adapter_001_src_channel;                                                                          // width_adapter_001:out_channel -> rsp_xbar_demux_004:sink_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                          // width_adapter_002:in_ready -> cmd_xbar_demux_004:src0_ready
	wire          width_adapter_002_src_endofpacket;                                                                      // width_adapter_002:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                            // width_adapter_002:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                    // width_adapter_002:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [75:0] width_adapter_002_src_data;                                                                             // width_adapter_002:out_data -> burst_adapter:sink0_data
	wire          width_adapter_002_src_ready;                                                                            // burst_adapter:sink0_ready -> width_adapter_002:out_ready
	wire    [1:0] width_adapter_002_src_channel;                                                                          // width_adapter_002:out_channel -> burst_adapter:sink0_channel
	wire          id_router_014_src_endofpacket;                                                                          // id_router_014:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_014_src_valid;                                                                                // id_router_014:src_valid -> width_adapter_003:in_valid
	wire          id_router_014_src_startofpacket;                                                                        // id_router_014:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [75:0] id_router_014_src_data;                                                                                 // id_router_014:src_data -> width_adapter_003:in_data
	wire    [1:0] id_router_014_src_channel;                                                                              // id_router_014:src_channel -> width_adapter_003:in_channel
	wire          id_router_014_src_ready;                                                                                // width_adapter_003:in_ready -> id_router_014:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                      // width_adapter_003:out_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                            // width_adapter_003:out_valid -> rsp_xbar_demux_014:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                    // width_adapter_003:out_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [93:0] width_adapter_003_src_data;                                                                             // width_adapter_003:out_data -> rsp_xbar_demux_014:sink_data
	wire          width_adapter_003_src_ready;                                                                            // rsp_xbar_demux_014:sink_ready -> width_adapter_003:out_ready
	wire    [1:0] width_adapter_003_src_channel;                                                                          // width_adapter_003:out_channel -> rsp_xbar_demux_014:sink_channel
	wire          crosser_out_endofpacket;                                                                                // crosser:out_endofpacket -> remote_update_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                      // crosser:out_valid -> remote_update_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                              // crosser:out_startofpacket -> remote_update_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] crosser_out_data;                                                                                       // crosser:out_data -> remote_update_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] crosser_out_channel;                                                                                    // crosser:out_channel -> remote_update_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src5_endofpacket;                                                                    // cmd_xbar_demux_003:src5_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_003_src5_valid;                                                                          // cmd_xbar_demux_003:src5_valid -> crosser:in_valid
	wire          cmd_xbar_demux_003_src5_startofpacket;                                                                  // cmd_xbar_demux_003:src5_startofpacket -> crosser:in_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src5_data;                                                                           // cmd_xbar_demux_003:src5_data -> crosser:in_data
	wire    [8:0] cmd_xbar_demux_003_src5_channel;                                                                        // cmd_xbar_demux_003:src5_channel -> crosser:in_channel
	wire          cmd_xbar_demux_003_src5_ready;                                                                          // crosser:in_ready -> cmd_xbar_demux_003:src5_ready
	wire          crosser_001_out_endofpacket;                                                                            // crosser_001:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_001_out_valid;                                                                                  // crosser_001:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_001_out_startofpacket;                                                                          // crosser_001:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] crosser_001_out_data;                                                                                   // crosser_001:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] crosser_001_out_channel;                                                                                // crosser_001:out_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src7_endofpacket;                                                                    // cmd_xbar_demux_003:src7_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_003_src7_valid;                                                                          // cmd_xbar_demux_003:src7_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_003_src7_startofpacket;                                                                  // cmd_xbar_demux_003:src7_startofpacket -> crosser_001:in_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src7_data;                                                                           // cmd_xbar_demux_003:src7_data -> crosser_001:in_data
	wire    [8:0] cmd_xbar_demux_003_src7_channel;                                                                        // cmd_xbar_demux_003:src7_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_003_src7_ready;                                                                          // crosser_001:in_ready -> cmd_xbar_demux_003:src7_ready
	wire          crosser_002_out_endofpacket;                                                                            // crosser_002:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_002_out_valid;                                                                                  // crosser_002:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_002_out_startofpacket;                                                                          // crosser_002:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] crosser_002_out_data;                                                                                   // crosser_002:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [8:0] crosser_002_out_channel;                                                                                // crosser_002:out_channel -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src8_endofpacket;                                                                    // cmd_xbar_demux_003:src8_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_003_src8_valid;                                                                          // cmd_xbar_demux_003:src8_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_003_src8_startofpacket;                                                                  // cmd_xbar_demux_003:src8_startofpacket -> crosser_002:in_startofpacket
	wire   [83:0] cmd_xbar_demux_003_src8_data;                                                                           // cmd_xbar_demux_003:src8_data -> crosser_002:in_data
	wire    [8:0] cmd_xbar_demux_003_src8_channel;                                                                        // cmd_xbar_demux_003:src8_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_003_src8_ready;                                                                          // crosser_002:in_ready -> cmd_xbar_demux_003:src8_ready
	wire          crosser_003_out_endofpacket;                                                                            // crosser_003:out_endofpacket -> rsp_xbar_mux_003:sink5_endofpacket
	wire          crosser_003_out_valid;                                                                                  // crosser_003:out_valid -> rsp_xbar_mux_003:sink5_valid
	wire          crosser_003_out_startofpacket;                                                                          // crosser_003:out_startofpacket -> rsp_xbar_mux_003:sink5_startofpacket
	wire   [83:0] crosser_003_out_data;                                                                                   // crosser_003:out_data -> rsp_xbar_mux_003:sink5_data
	wire    [8:0] crosser_003_out_channel;                                                                                // crosser_003:out_channel -> rsp_xbar_mux_003:sink5_channel
	wire          crosser_003_out_ready;                                                                                  // rsp_xbar_mux_003:sink5_ready -> crosser_003:out_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                    // rsp_xbar_demux_010:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                          // rsp_xbar_demux_010:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                  // rsp_xbar_demux_010:src0_startofpacket -> crosser_003:in_startofpacket
	wire   [83:0] rsp_xbar_demux_010_src0_data;                                                                           // rsp_xbar_demux_010:src0_data -> crosser_003:in_data
	wire    [8:0] rsp_xbar_demux_010_src0_channel;                                                                        // rsp_xbar_demux_010:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                          // crosser_003:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          crosser_004_out_endofpacket;                                                                            // crosser_004:out_endofpacket -> rsp_xbar_mux_003:sink7_endofpacket
	wire          crosser_004_out_valid;                                                                                  // crosser_004:out_valid -> rsp_xbar_mux_003:sink7_valid
	wire          crosser_004_out_startofpacket;                                                                          // crosser_004:out_startofpacket -> rsp_xbar_mux_003:sink7_startofpacket
	wire   [83:0] crosser_004_out_data;                                                                                   // crosser_004:out_data -> rsp_xbar_mux_003:sink7_data
	wire    [8:0] crosser_004_out_channel;                                                                                // crosser_004:out_channel -> rsp_xbar_mux_003:sink7_channel
	wire          crosser_004_out_ready;                                                                                  // rsp_xbar_mux_003:sink7_ready -> crosser_004:out_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                    // rsp_xbar_demux_012:src0_endofpacket -> crosser_004:in_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                          // rsp_xbar_demux_012:src0_valid -> crosser_004:in_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                  // rsp_xbar_demux_012:src0_startofpacket -> crosser_004:in_startofpacket
	wire   [83:0] rsp_xbar_demux_012_src0_data;                                                                           // rsp_xbar_demux_012:src0_data -> crosser_004:in_data
	wire    [8:0] rsp_xbar_demux_012_src0_channel;                                                                        // rsp_xbar_demux_012:src0_channel -> crosser_004:in_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                          // crosser_004:in_ready -> rsp_xbar_demux_012:src0_ready
	wire          crosser_005_out_endofpacket;                                                                            // crosser_005:out_endofpacket -> rsp_xbar_mux_003:sink8_endofpacket
	wire          crosser_005_out_valid;                                                                                  // crosser_005:out_valid -> rsp_xbar_mux_003:sink8_valid
	wire          crosser_005_out_startofpacket;                                                                          // crosser_005:out_startofpacket -> rsp_xbar_mux_003:sink8_startofpacket
	wire   [83:0] crosser_005_out_data;                                                                                   // crosser_005:out_data -> rsp_xbar_mux_003:sink8_data
	wire    [8:0] crosser_005_out_channel;                                                                                // crosser_005:out_channel -> rsp_xbar_mux_003:sink8_channel
	wire          crosser_005_out_ready;                                                                                  // rsp_xbar_mux_003:sink8_ready -> crosser_005:out_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                    // rsp_xbar_demux_013:src0_endofpacket -> crosser_005:in_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                          // rsp_xbar_demux_013:src0_valid -> crosser_005:in_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                  // rsp_xbar_demux_013:src0_startofpacket -> crosser_005:in_startofpacket
	wire   [83:0] rsp_xbar_demux_013_src0_data;                                                                           // rsp_xbar_demux_013:src0_data -> crosser_005:in_data
	wire    [8:0] rsp_xbar_demux_013_src0_channel;                                                                        // rsp_xbar_demux_013:src0_channel -> crosser_005:in_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                          // crosser_005:in_ready -> rsp_xbar_demux_013:src0_ready
	wire    [3:0] limiter_cmd_valid_data;                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [3:0] limiter_001_cmd_valid_data;                                                                             // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire    [8:0] limiter_002_cmd_valid_data;                                                                             // limiter_002:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire    [1:0] limiter_003_cmd_valid_data;                                                                             // limiter_003:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire   [31:0] cpu_d_irq_irq;                                                                                          // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver0_irq;                                                                               // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                          // button_pio:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                                                               // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                      // high_res_timer:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                               // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                      // jtag_uart:av_irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver3_irq;                                                                               // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                                      // sys_clk_timer:irq -> irq_synchronizer_003:receiver_irq

	cycloneIII_3c25_niosII_standard_sopc_ddr_sdram ddr_sdram (
		.local_address     (ddr_sdram_s1_translator_avalon_anti_slave_0_address),            //                  s1.address
		.local_write_req   (ddr_sdram_s1_translator_avalon_anti_slave_0_write),              //                    .write
		.local_read_req    (ddr_sdram_s1_translator_avalon_anti_slave_0_read),               //                    .read
		.local_burstbegin  (ddr_sdram_s1_translator_avalon_anti_slave_0_beginbursttransfer), //                    .beginbursttransfer
		.local_ready       (ddr_sdram_s1_translator_avalon_anti_slave_0_waitrequest),        //                    .waitrequest_n
		.local_rdata       (ddr_sdram_s1_translator_avalon_anti_slave_0_readdata),           //                    .readdata
		.local_rdata_valid (ddr_sdram_s1_translator_avalon_anti_slave_0_readdatavalid),      //                    .readdatavalid
		.local_wdata       (ddr_sdram_s1_translator_avalon_anti_slave_0_writedata),          //                    .writedata
		.local_be          (ddr_sdram_s1_translator_avalon_anti_slave_0_byteenable),         //                    .byteenable
		.local_size        (ddr_sdram_s1_translator_avalon_anti_slave_0_burstcount),         //                    .burstcount
		.local_refresh_ack (local_refresh_ack_from_the_ddr_sdram),                           // external_connection.export
		.local_wdata_req   (local_wdata_req_from_the_ddr_sdram),                             //                    .export
		.local_init_done   (local_init_done_from_the_ddr_sdram),                             //                    .export
		.reset_phy_clk_n   (reset_phy_clk_n_from_the_ddr_sdram),                             //                    .export
		.mem_clk           (mem_clk_to_and_from_the_ddr_sdram),                              //              memory.mem_clk
		.mem_clk_n         (mem_clk_n_to_and_from_the_ddr_sdram),                            //                    .mem_clk_n
		.mem_cs_n          (mem_cs_n_from_the_ddr_sdram),                                    //                    .mem_cs_n
		.mem_cke           (mem_cke_from_the_ddr_sdram),                                     //                    .mem_cke
		.mem_addr          (mem_addr_from_the_ddr_sdram),                                    //                    .mem_addr
		.mem_ba            (mem_ba_from_the_ddr_sdram),                                      //                    .mem_ba
		.mem_ras_n         (mem_ras_n_from_the_ddr_sdram),                                   //                    .mem_ras_n
		.mem_cas_n         (mem_cas_n_from_the_ddr_sdram),                                   //                    .mem_cas_n
		.mem_we_n          (mem_we_n_from_the_ddr_sdram),                                    //                    .mem_we_n
		.mem_dq            (mem_dq_to_and_from_the_ddr_sdram),                               //                    .mem_dq
		.mem_dqs           (mem_dqs_to_and_from_the_ddr_sdram),                              //                    .mem_dqs
		.mem_dm            (mem_dm_from_the_ddr_sdram),                                      //                    .mem_dm
		.pll_ref_clk       (clk),                                                            //              refclk.clk
		.soft_reset_n      (~rst_controller_reset_out_reset),                                //        soft_reset_n.reset_n
		.global_reset_n    (ddr_sdram_reset_n),                                              //      global_reset_n.reset_n
		.reset_request_n   (ddr_sdram_reset_request_n_reset),                                //     reset_request_n.reset_n
		.phy_clk           (ddr_sdram_phy_clk_out),                                          //              sysclk.clk
		.aux_full_rate_clk (ddr_sdram_aux_full_rate_clk_out),                                //             auxfull.clk
		.aux_half_rate_clk (ddr_sdram_aux_half_rate_clk_out)                                 //             auxhalf.clk
	);

	cycloneIII_3c25_niosII_standard_sopc_sys_clk_timer sys_clk_timer (
		.clk        (pll_c2_out),                                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_003_receiver_irq)                           //   irq.irq
	);

	cycloneIII_3c25_niosII_standard_sopc_high_res_timer high_res_timer (
		.clk        (pll_c2_out),                                                  //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         // reset.reset_n
		.address    (high_res_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_res_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                            //   irq.irq
	);

	cycloneIII_3c25_niosII_standard_sopc_performance_counter performance_counter (
		.clk           (pll_c2_out),                                                                     //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                                            //         reset.reset_n
		.address       (performance_counter_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	cycloneIII_3c25_niosII_standard_sopc_jtag_uart jtag_uart (
		.clk            (pll_c2_out),                                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_002_receiver_irq)                                       //               irq.irq
	);

	cycloneIII_3c25_niosII_standard_sopc_button_pio button_pio (
		.clk        (pll_c2_out),                                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (in_port_to_the_button_pio),                               // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)                            //                 irq.irq
	);

	cycloneIII_3c25_niosII_standard_sopc_led_pio led_pio (
		.clk        (pll_c2_out),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led_pio)                             // external_connection.export
	);

	altera_avalon_remote_update_cycloneiii remote_update (
		.clk         (pll_c3_out),                                                  //       global_signals_clock.clk
		.reset       (rst_controller_002_reset_out_reset),                          // global_signals_clock_reset.reset
		.writedata   (remote_update_s1_translator_avalon_anti_slave_0_writedata),   //                         s1.writedata
		.readdata    (remote_update_s1_translator_avalon_anti_slave_0_readdata),    //                           .readdata
		.address     (remote_update_s1_translator_avalon_anti_slave_0_address),     //                           .address
		.chipselect  (remote_update_s1_translator_avalon_anti_slave_0_chipselect),  //                           .chipselect
		.write       (remote_update_s1_translator_avalon_anti_slave_0_write),       //                           .write
		.read        (remote_update_s1_translator_avalon_anti_slave_0_read),        //                           .read
		.waitrequest (remote_update_s1_translator_avalon_anti_slave_0_waitrequest)  //                           .waitrequest
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (25),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) flash_ssram_pipeline_bridge (
		.clk              (pll_c0_out),                                                                  //   clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                          // reset.reset
		.s0_waitrequest   (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (flash_ssram_pipeline_bridge_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (flash_ssram_pipeline_bridge_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (flash_ssram_pipeline_bridge_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (flash_ssram_pipeline_bridge_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (flash_ssram_pipeline_bridge_m0_writedata),                                    //      .writedata
		.m0_address       (flash_ssram_pipeline_bridge_m0_address),                                      //      .address
		.m0_write         (flash_ssram_pipeline_bridge_m0_write),                                        //      .write
		.m0_read          (flash_ssram_pipeline_bridge_m0_read),                                         //      .read
		.m0_byteenable    (flash_ssram_pipeline_bridge_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (flash_ssram_pipeline_bridge_m0_debugaccess)                                   //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (25),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipeline_bridge_before_tristate_bridge (
		.clk              (pll_c0_out),                                              //   clk.clk
		.reset            (rst_controller_003_reset_out_reset),                      // reset.reset
		.s0_waitrequest   (flash_ssram_pipeline_bridge_m0_waitrequest),              //    s0.waitrequest
		.s0_readdata      (flash_ssram_pipeline_bridge_m0_readdata),                 //      .readdata
		.s0_readdatavalid (flash_ssram_pipeline_bridge_m0_readdatavalid),            //      .readdatavalid
		.s0_burstcount    (flash_ssram_pipeline_bridge_m0_burstcount),               //      .burstcount
		.s0_writedata     (flash_ssram_pipeline_bridge_m0_writedata),                //      .writedata
		.s0_address       (flash_ssram_pipeline_bridge_m0_address),                  //      .address
		.s0_write         (flash_ssram_pipeline_bridge_m0_write),                    //      .write
		.s0_read          (flash_ssram_pipeline_bridge_m0_read),                     //      .read
		.s0_byteenable    (flash_ssram_pipeline_bridge_m0_byteenable),               //      .byteenable
		.s0_debugaccess   (flash_ssram_pipeline_bridge_m0_debugaccess),              //      .debugaccess
		.m0_waitrequest   (pipeline_bridge_before_tristate_bridge_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (pipeline_bridge_before_tristate_bridge_m0_readdata),      //      .readdata
		.m0_readdatavalid (pipeline_bridge_before_tristate_bridge_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (pipeline_bridge_before_tristate_bridge_m0_burstcount),    //      .burstcount
		.m0_writedata     (pipeline_bridge_before_tristate_bridge_m0_writedata),     //      .writedata
		.m0_address       (pipeline_bridge_before_tristate_bridge_m0_address),       //      .address
		.m0_write         (pipeline_bridge_before_tristate_bridge_m0_write),         //      .write
		.m0_read          (pipeline_bridge_before_tristate_bridge_m0_read),          //      .read
		.m0_byteenable    (pipeline_bridge_before_tristate_bridge_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (pipeline_bridge_before_tristate_bridge_m0_debugaccess)    //      .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (25),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_ddr_clock_bridge (
		.m0_clk           (ddr_sdram_phy_clk_out),                                                //   m0_clk.clk
		.m0_reset         (rst_controller_004_reset_out_reset),                                   // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                           //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                                   // s0_reset.reset
		.s0_waitrequest   (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_ddr_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (cpu_ddr_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (cpu_ddr_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (cpu_ddr_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (cpu_ddr_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (cpu_ddr_clock_bridge_m0_address),                                      //         .address
		.m0_write         (cpu_ddr_clock_bridge_m0_write),                                        //         .write
		.m0_read          (cpu_ddr_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (cpu_ddr_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (cpu_ddr_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) slow_peripheral_bridge (
		.m0_clk           (pll_c2_out),                                                             //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                                     // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                             //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                                     // s0_reset.reset
		.s0_waitrequest   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_peripheral_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (slow_peripheral_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (slow_peripheral_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (slow_peripheral_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (slow_peripheral_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (slow_peripheral_bridge_m0_address),                                      //         .address
		.m0_write         (slow_peripheral_bridge_m0_write),                                        //         .write
		.m0_read          (slow_peripheral_bridge_m0_read),                                         //         .read
		.m0_byteenable    (slow_peripheral_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (slow_peripheral_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	cycloneIII_3c25_niosII_standard_sopc_cpu cpu (
		.clk                                   (pll_c0_out),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_003_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	cycloneIII_3c25_niosII_standard_sopc_sysid sysid (
		.clock    (pll_c0_out),                                                  //           clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	cycloneIII_3c25_niosII_standard_sopc_flash_ssram_tristate_bridge_bridge_0 flash_ssram_tristate_bridge_bridge_0 (
		.clk                                        (pll_c0_out),                                                                          //   clk.clk
		.reset                                      (rst_controller_003_reset_out_reset),                                                  // reset.reset
		.request                                    (flash_ssram_tristate_bridge_pinsharer_0_tcm_request),                                 //   tcs.request
		.grant                                      (flash_ssram_tristate_bridge_pinsharer_0_tcm_grant),                                   //      .grant
		.tcs_read_n_to_the_ext_flash                (flash_ssram_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out),             //      .read_n_to_the_ext_flash_out
		.tcs_select_n_to_the_ext_flash              (flash_ssram_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),           //      .select_n_to_the_ext_flash_out
		.tcs_flash_ssram_tristate_bridge_address    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_address_out), //      .flash_ssram_tristate_bridge_address_out
		.tcs_bwe_n_to_the_ssram                     (flash_ssram_tristate_bridge_pinsharer_0_tcm_bwe_n_to_the_ssram_out),                  //      .bwe_n_to_the_ssram_out
		.tcs_reset_n_to_the_ssram                   (flash_ssram_tristate_bridge_pinsharer_0_tcm_reset_n_to_the_ssram_out),                //      .reset_n_to_the_ssram_out
		.tcs_chipenable1_n_to_the_ssram             (flash_ssram_tristate_bridge_pinsharer_0_tcm_chipenable1_n_to_the_ssram_out),          //      .chipenable1_n_to_the_ssram_out
		.tcs_bw_n_to_the_ssram                      (flash_ssram_tristate_bridge_pinsharer_0_tcm_bw_n_to_the_ssram_out),                   //      .bw_n_to_the_ssram_out
		.tcs_outputenable_n_to_the_ssram            (flash_ssram_tristate_bridge_pinsharer_0_tcm_outputenable_n_to_the_ssram_out),         //      .outputenable_n_to_the_ssram_out
		.tcs_flash_ssram_tristate_bridge_data       (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_out),    //      .flash_ssram_tristate_bridge_data_out
		.tcs_flash_ssram_tristate_bridge_data_outen (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_outen),  //      .flash_ssram_tristate_bridge_data_outen
		.tcs_flash_ssram_tristate_bridge_data_in    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_in),     //      .flash_ssram_tristate_bridge_data_in
		.tcs_adsc_n_to_the_ssram                    (flash_ssram_tristate_bridge_pinsharer_0_tcm_adsc_n_to_the_ssram_out),                 //      .adsc_n_to_the_ssram_out
		.tcs_write_n_to_the_ext_flash               (flash_ssram_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out),            //      .write_n_to_the_ext_flash_out
		.read_n_to_the_ext_flash                    (read_n_to_the_ext_flash),                                                             //   out.read_n_to_the_ext_flash
		.select_n_to_the_ext_flash                  (select_n_to_the_ext_flash),                                                           //      .select_n_to_the_ext_flash
		.flash_ssram_tristate_bridge_address        (flash_ssram_tristate_bridge_address),                                                 //      .flash_ssram_tristate_bridge_address
		.bwe_n_to_the_ssram                         (bwe_n_to_the_ssram),                                                                  //      .bwe_n_to_the_ssram
		.reset_n_to_the_ssram                       (reset_n_to_the_ssram),                                                                //      .reset_n_to_the_ssram
		.chipenable1_n_to_the_ssram                 (chipenable1_n_to_the_ssram),                                                          //      .chipenable1_n_to_the_ssram
		.bw_n_to_the_ssram                          (bw_n_to_the_ssram),                                                                   //      .bw_n_to_the_ssram
		.outputenable_n_to_the_ssram                (outputenable_n_to_the_ssram),                                                         //      .outputenable_n_to_the_ssram
		.flash_ssram_tristate_bridge_data           (flash_ssram_tristate_bridge_data),                                                    //      .flash_ssram_tristate_bridge_data
		.adsc_n_to_the_ssram                        (adsc_n_to_the_ssram),                                                                 //      .adsc_n_to_the_ssram
		.write_n_to_the_ext_flash                   (write_n_to_the_ext_flash)                                                             //      .write_n_to_the_ext_flash
	);

	cycloneIII_3c25_niosII_standard_sopc_flash_ssram_tristate_bridge_pinSharer_0 flash_ssram_tristate_bridge_pinsharer_0 (
		.clk_clk                                (pll_c0_out),                                                                          //   clk.clk
		.reset_reset                            (rst_controller_003_reset_out_reset),                                                  // reset.reset
		.request                                (flash_ssram_tristate_bridge_pinsharer_0_tcm_request),                                 //   tcm.request
		.grant                                  (flash_ssram_tristate_bridge_pinsharer_0_tcm_grant),                                   //      .grant
		.chipenable1_n_to_the_ssram             (flash_ssram_tristate_bridge_pinsharer_0_tcm_chipenable1_n_to_the_ssram_out),          //      .chipenable1_n_to_the_ssram_out
		.bw_n_to_the_ssram                      (flash_ssram_tristate_bridge_pinsharer_0_tcm_bw_n_to_the_ssram_out),                   //      .bw_n_to_the_ssram_out
		.outputenable_n_to_the_ssram            (flash_ssram_tristate_bridge_pinsharer_0_tcm_outputenable_n_to_the_ssram_out),         //      .outputenable_n_to_the_ssram_out
		.bwe_n_to_the_ssram                     (flash_ssram_tristate_bridge_pinsharer_0_tcm_bwe_n_to_the_ssram_out),                  //      .bwe_n_to_the_ssram_out
		.reset_n_to_the_ssram                   (flash_ssram_tristate_bridge_pinsharer_0_tcm_reset_n_to_the_ssram_out),                //      .reset_n_to_the_ssram_out
		.adsc_n_to_the_ssram                    (flash_ssram_tristate_bridge_pinsharer_0_tcm_adsc_n_to_the_ssram_out),                 //      .adsc_n_to_the_ssram_out
		.flash_ssram_tristate_bridge_address    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_address_out), //      .flash_ssram_tristate_bridge_address_out
		.read_n_to_the_ext_flash                (flash_ssram_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out),             //      .read_n_to_the_ext_flash_out
		.write_n_to_the_ext_flash               (flash_ssram_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out),            //      .write_n_to_the_ext_flash_out
		.flash_ssram_tristate_bridge_data       (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_out),    //      .flash_ssram_tristate_bridge_data_out
		.flash_ssram_tristate_bridge_data_in    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_in),     //      .flash_ssram_tristate_bridge_data_in
		.flash_ssram_tristate_bridge_data_outen (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_outen),  //      .flash_ssram_tristate_bridge_data_outen
		.select_n_to_the_ext_flash              (flash_ssram_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),           //      .select_n_to_the_ext_flash_out
		.tcs0_request                           (ext_flash_tcm_request),                                                               //  tcs0.request
		.tcs0_grant                             (ext_flash_tcm_grant),                                                                 //      .grant
		.tcs0_address_out                       (ext_flash_tcm_address_out),                                                           //      .address_out
		.tcs0_read_n_out                        (ext_flash_tcm_read_n_out),                                                            //      .read_n_out
		.tcs0_write_n_out                       (ext_flash_tcm_write_n_out),                                                           //      .write_n_out
		.tcs0_data_out                          (ext_flash_tcm_data_out),                                                              //      .data_out
		.tcs0_data_in                           (ext_flash_tcm_data_in),                                                               //      .data_in
		.tcs0_data_outen                        (ext_flash_tcm_data_outen),                                                            //      .data_outen
		.tcs0_chipselect_n_out                  (ext_flash_tcm_chipselect_n_out),                                                      //      .chipselect_n_out
		.tcs1_request                           (ssram_tcm_request),                                                                   //  tcs1.request
		.tcs1_grant                             (ssram_tcm_grant),                                                                     //      .grant
		.tcs1_chipselect_n_out                  (ssram_tcm_chipselect_n_out),                                                          //      .chipselect_n_out
		.tcs1_byteenable_n_out                  (ssram_tcm_byteenable_n_out),                                                          //      .byteenable_n_out
		.tcs1_outputenable_n_out                (ssram_tcm_outputenable_n_out),                                                        //      .outputenable_n_out
		.tcs1_write_n_out                       (ssram_tcm_write_n_out),                                                               //      .write_n_out
		.tcs1_data_out                          (ssram_tcm_data_out),                                                                  //      .data_out
		.tcs1_data_in                           (ssram_tcm_data_in),                                                                   //      .data_in
		.tcs1_data_outen                        (ssram_tcm_data_outen),                                                                //      .data_outen
		.tcs1_address_out                       (ssram_tcm_address_out),                                                               //      .address_out
		.tcs1_reset_n_out                       (ssram_tcm_reset_n_out),                                                               //      .reset_n_out
		.tcs1_begintransfer_n_out               (ssram_tcm_begintransfer_n_out)                                                        //      .begintransfer_n_out
	);

	cycloneIII_3c25_niosII_standard_sopc_ext_flash #(
		.TCM_ADDRESS_W                  (24),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (100),
		.TCM_WRITE_WAIT                 (100),
		.TCM_SETUP_WAIT                 (25),
		.TCM_DATA_HOLD                  (20),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash (
		.clk_clk              (pll_c0_out),                                                 //   clk.clk
		.reset_reset          (rst_controller_003_reset_out_reset),                         // reset.reset
		.uas_address          (ext_flash_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (ext_flash_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (ext_flash_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (ext_flash_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (ext_flash_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (ext_flash_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                                      //      .request
		.tcm_grant            (ext_flash_tcm_grant),                                        //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                                       //      .data_in
	);

	cycloneIII_3c25_niosII_standard_sopc_ssram #(
		.TCM_ADDRESS_W                  (20),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (0),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (1),
		.TCM_READLATENCY                (4),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (1),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (1),
		.CHIPSELECT_THROUGH_READLATENCY (1)
	) ssram (
		.clk_clk                 (pll_c0_out),                                             //   clk.clk
		.reset_reset             (rst_controller_003_reset_out_reset),                     // reset.reset
		.uas_address             (ssram_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount          (ssram_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read                (ssram_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write               (ssram_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest         (ssram_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid       (ssram_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable          (ssram_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata            (ssram_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata           (ssram_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock                (ssram_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess         (ssram_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out         (ssram_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_begintransfer_n_out (ssram_tcm_begintransfer_n_out),                          //      .begintransfer_n_out
		.tcm_chipselect_n_out    (ssram_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_outputenable_n_out  (ssram_tcm_outputenable_n_out),                           //      .outputenable_n_out
		.tcm_reset_n_out         (ssram_tcm_reset_n_out),                                  //      .reset_n_out
		.tcm_request             (ssram_tcm_request),                                      //      .request
		.tcm_grant               (ssram_tcm_grant),                                        //      .grant
		.tcm_address_out         (ssram_tcm_address_out),                                  //      .address_out
		.tcm_byteenable_n_out    (ssram_tcm_byteenable_n_out),                             //      .byteenable_n_out
		.tcm_data_out            (ssram_tcm_data_out),                                     //      .data_out
		.tcm_data_outen          (ssram_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in             (ssram_tcm_data_in)                                       //      .data_in
	);

	cycloneIII_3c25_niosII_standard_sopc_pll pll (
		.clk       (clk),                                                    //       inclk_interface.clk
		.reset     (rst_controller_005_reset_out_reset),                     // inclk_interface_reset.reset
		.read      (pll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (pll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (pll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (pll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (pll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (pll_c0_out),                                             //                    c0.clk
		.c1        (pll_c1_clk),                                             //                    c1.clk
		.c2        (pll_c2_out),                                             //                    c2.clk
		.c3        (pll_c3_out),                                             //                    c3.clk
		.areset    (pll_areset_conduit_export),                              //        areset_conduit.export
		.locked    (pll_locked_conduit_export),                              //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)                            //     phasedone_conduit.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (pll_c0_out),                                                         //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                 //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (28),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (pll_c0_out),                                                                //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                        //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (pll_c0_out),                                                                       //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                               //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) flash_ssram_pipeline_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                                //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                        //                    reset.reset
		.uav_address           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_chipselect         (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_ddr_clock_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                         //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (28),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slow_peripheral_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                           //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_ddr_clock_bridge_m0_translator (
		.clk                   (ddr_sdram_phy_clk_out),                                                      //                       clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                         //                     reset.reset
		.uav_address           (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_ddr_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_ddr_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (cpu_ddr_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (cpu_ddr_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (cpu_ddr_clock_bridge_m0_read),                                               //                          .read
		.av_readdata           (cpu_ddr_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_ddr_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_ddr_clock_bridge_m0_write),                                              //                          .write
		.av_writedata          (cpu_ddr_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_ddr_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                       //               (terminated)
		.av_begintransfer      (1'b0),                                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                                       //               (terminated)
		.av_lock               (1'b0),                                                                       //               (terminated)
		.uav_clken             (),                                                                           //               (terminated)
		.av_clken              (1'b1)                                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr_sdram_s1_translator (
		.clk                   (ddr_sdram_phy_clk_out),                                                   //                      clk.clk
		.reset                 (~ddr_sdram_reset_request_n_reset),                                        //                    reset.reset
		.uav_address           (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ddr_sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ddr_sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ddr_sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ddr_sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ddr_sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer (ddr_sdram_s1_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount         (ddr_sdram_s1_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ddr_sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ddr_sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (~ddr_sdram_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_chipselect         (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (9),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (9),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) slow_peripheral_bridge_m0_translator (
		.clk                   (pll_c2_out),                                                                   //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (slow_peripheral_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (slow_peripheral_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (slow_peripheral_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (slow_peripheral_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (slow_peripheral_bridge_m0_read),                                               //                          .read
		.av_readdata           (slow_peripheral_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (slow_peripheral_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (slow_peripheral_bridge_m0_write),                                              //                          .write
		.av_writedata          (slow_peripheral_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (slow_peripheral_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                   (pll_c2_out),                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_res_timer_s1_translator (
		.clk                   (pll_c2_out),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_res_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_res_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (pll_c2_out),                                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_pio_s1_translator (
		.clk                   (pll_c2_out),                                                            //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_control_slave_translator (
		.clk                   (pll_c2_out),                                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (performance_counter_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (performance_counter_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read               (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_byteenable         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_chipselect         (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (6),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (2),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) remote_update_s1_translator (
		.clk                   (pll_c3_out),                                                                  //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                          //                    reset.reset
		.uav_address           (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (remote_update_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (remote_update_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (remote_update_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (remote_update_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (remote_update_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (remote_update_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (remote_update_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                   (pll_c2_out),                                                                  //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (pll_c0_out),                                                                     //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                             //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (9),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pll_pll_slave_translator (
		.clk                   (clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                       //                    reset.reset
		.uav_address           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pipeline_bridge_before_tristate_bridge_m0_translator (
		.clk                   (pll_c0_out),                                                                                   //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                           //                     reset.reset
		.uav_address           (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (pipeline_bridge_before_tristate_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (pipeline_bridge_before_tristate_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (pipeline_bridge_before_tristate_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (pipeline_bridge_before_tristate_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (pipeline_bridge_before_tristate_bridge_m0_read),                                               //                          .read
		.av_readdata           (pipeline_bridge_before_tristate_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (pipeline_bridge_before_tristate_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (pipeline_bridge_before_tristate_bridge_m0_write),                                              //                          .write
		.av_writedata          (pipeline_bridge_before_tristate_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (pipeline_bridge_before_tristate_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                                         //               (terminated)
		.uav_clken             (),                                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (2),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ext_flash_uas_translator (
		.clk                   (pll_c0_out),                                                               //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                       //                    reset.reset
		.uav_address           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ext_flash_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ext_flash_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ext_flash_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ext_flash_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ext_flash_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (ext_flash_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ssram_uas_translator (
		.clk                   (pll_c0_out),                                                           //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                   //                    reset.reset
		.uav_address           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ssram_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ssram_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ssram_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ssram_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ssram_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ssram_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (ssram_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ssram_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ssram_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (ssram_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (ssram_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (ssram_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                  //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                          // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                        //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                        //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (83),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_TRANS_EXCLUSIVE       (69),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (82),
		.PKT_DATA_SIDEBAND_L       (82),
		.PKT_QOS_H                 (84),
		.PKT_QOS_L                 (84),
		.PKT_ADDR_SIDEBAND_H       (81),
		.PKT_ADDR_SIDEBAND_L       (81),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                         //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                           //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                 //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                 //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                          //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                        //                .channel
		.rf_sink_ready           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (11),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                   //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                 //                .channel
		.rf_sink_ready           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                   //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (63),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (64),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.PKT_TRANS_READ            (67),
		.PKT_TRANS_LOCK            (68),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                     //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                                    //                .channel
		.rf_sink_ready           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (81),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                     //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_BEGIN_BURST           (82),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.PKT_BURST_TYPE_H          (79),
		.PKT_BURST_TYPE_L          (78),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (86),
		.PKT_THREAD_ID_L           (86),
		.PKT_CACHE_H               (93),
		.PKT_CACHE_L               (90),
		.PKT_DATA_SIDEBAND_H       (81),
		.PKT_DATA_SIDEBAND_L       (81),
		.PKT_QOS_H                 (83),
		.PKT_QOS_L                 (83),
		.PKT_ADDR_SIDEBAND_H       (80),
		.PKT_ADDR_SIDEBAND_L       (80),
		.ST_DATA_W                 (96),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (15),
		.CACHE_VALUE               (4'b0000)
	) cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (ddr_sdram_phy_clk_out),                                                               //       clk.clk
		.reset            (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_004_src0_valid),                                                       //        rp.valid
		.rp_data          (rsp_xbar_demux_004_src0_data),                                                        //          .data
		.rp_channel       (rsp_xbar_demux_004_src0_channel),                                                     //          .channel
		.rp_startofpacket (rsp_xbar_demux_004_src0_startofpacket),                                               //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),                                                 //          .endofpacket
		.rp_ready         (rsp_xbar_demux_004_src0_ready)                                                        //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (118),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (96),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (97),
		.PKT_TRANS_POSTED          (98),
		.PKT_TRANS_WRITE           (99),
		.PKT_TRANS_READ            (100),
		.PKT_TRANS_LOCK            (101),
		.PKT_SRC_ID_H              (120),
		.PKT_SRC_ID_L              (120),
		.PKT_DEST_ID_H             (121),
		.PKT_DEST_ID_L             (121),
		.PKT_BURSTWRAP_H           (110),
		.PKT_BURSTWRAP_L           (107),
		.PKT_BYTE_CNT_H            (106),
		.PKT_BYTE_CNT_L            (103),
		.PKT_PROTECTION_H          (125),
		.PKT_PROTECTION_L          (123),
		.PKT_RESPONSE_STATUS_H     (131),
		.PKT_RESPONSE_STATUS_L     (130),
		.PKT_BURST_SIZE_H          (113),
		.PKT_BURST_SIZE_L          (111),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (132),
		.AVS_BURSTCOUNT_W          (4),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ddr_sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr_sdram_phy_clk_out),                                                             //             clk.clk
		.reset                   (~ddr_sdram_reset_request_n_reset),                                                  //       clk_reset.reset
		.m0_address              (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (width_adapter_src_ready),                                                           //              cp.ready
		.cp_valid                (width_adapter_src_valid),                                                           //                .valid
		.cp_data                 (width_adapter_src_data),                                                            //                .data
		.cp_startofpacket        (width_adapter_src_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (width_adapter_src_endofpacket),                                                     //                .endofpacket
		.cp_channel              (width_adapter_src_channel),                                                         //                .channel
		.rf_sink_ready           (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (133),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr_sdram_phy_clk_out),                                                             //       clk.clk
		.reset             (~ddr_sdram_reset_request_n_reset),                                                  // clk_reset.reset
		.in_data           (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (64),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.PKT_BURST_TYPE_H          (61),
		.PKT_BURST_TYPE_L          (60),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_TRANS_EXCLUSIVE       (50),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_DATA_SIDEBAND_H       (63),
		.PKT_DATA_SIDEBAND_L       (63),
		.PKT_QOS_H                 (65),
		.PKT_QOS_L                 (65),
		.PKT_ADDR_SIDEBAND_H       (62),
		.PKT_ADDR_SIDEBAND_L       (62),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (pll_c2_out),                                                                            //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src0_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src0_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_003_src0_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src0_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src0_channel),                                                    //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src1_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src1_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_003_src1_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src1_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src1_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src1_channel),                                                        //                .channel
		.rf_sink_ready           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_003_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src3_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src3_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_003_src3_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src3_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src3_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src3_channel),                                                 //                .channel
		.rf_sink_ready           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src4_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src4_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_003_src4_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src4_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src4_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src4_channel),                                                                        //                .channel
		.rf_sink_ready           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) remote_update_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (remote_update_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                     //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                     //                .valid
		.cp_data                 (crosser_out_data),                                                                      //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                               //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                   //                .channel
		.rf_sink_ready           (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (remote_update_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (remote_update_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c3_out),                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (remote_update_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src6_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src6_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_003_src6_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src6_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src6_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src6_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                               //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                    //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                    //                .valid
		.cp_data                 (crosser_001_out_data),                                                                     //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                              //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                  //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                              //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                              //                .valid
		.cp_data                 (crosser_002_out_data),                                                               //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                        //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                            //                .channel
		.rf_sink_ready           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk),                                                                          //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                           // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (83),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                                            //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                                    // clk_reset.reset
		.av_address       (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_003_rsp_src_valid),                                                                             //        rp.valid
		.rp_data          (limiter_003_rsp_src_data),                                                                              //          .data
		.rp_channel       (limiter_003_rsp_src_channel),                                                                           //          .channel
		.rp_startofpacket (limiter_003_rsp_src_startofpacket),                                                                     //          .startofpacket
		.rp_endofpacket   (limiter_003_rsp_src_endofpacket),                                                                       //          .endofpacket
		.rp_ready         (limiter_003_rsp_src_ready)                                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (65),
		.PKT_DEST_ID_L             (65),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (69),
		.PKT_PROTECTION_L          (67),
		.PKT_RESPONSE_STATUS_H     (75),
		.PKT_RESPONSE_STATUS_L     (74),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                         //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ssram_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                     //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ssram_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ssram_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_004_src1_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_004_src1_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_004_src1_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_004_src1_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_004_src1_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_004_src1_channel),                                                //                .channel
		.rf_sink_ready           (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (6),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                     //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.in_data           (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	cycloneIII_3c25_niosII_standard_sopc_addr_router addr_router (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                       //          .valid
		.src_data           (addr_router_src_data),                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                  //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router id_router_001 (
		.sink_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                              //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router id_router_002 (
		.sink_ready         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                            //       src.ready
		.src_valid          (id_router_002_src_valid),                                                            //          .valid
		.src_data           (id_router_002_src_data),                                                             //          .data
		.src_channel        (id_router_002_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                       //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_003 id_router_003 (
		.sink_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                           //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                              //       src.ready
		.src_valid          (id_router_003_src_valid),                                                              //          .valid
		.src_data           (id_router_003_src_data),                                                               //          .data
		.src_channel        (id_router_003_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                         //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_addr_router_002 addr_router_002 (
		.sink_ready         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr_sdram_phy_clk_out),                                                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                           //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                           //          .valid
		.src_data           (addr_router_002_src_data),                                                            //          .data
		.src_channel        (addr_router_002_src_channel),                                                         //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                      //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_004 id_router_004 (
		.sink_ready         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr_sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr_sdram_phy_clk_out),                                                   //       clk.clk
		.reset              (~ddr_sdram_reset_request_n_reset),                                        // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                 //       src.ready
		.src_valid          (id_router_004_src_valid),                                                 //          .valid
		.src_data           (id_router_004_src_data),                                                  //          .data
		.src_channel        (id_router_004_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                            //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_addr_router_003 addr_router_003 (
		.sink_ready         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_005 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                  //       src.ready
		.src_valid          (id_router_005_src_valid),                                                  //          .valid
		.src_data           (id_router_005_src_data),                                                   //          .data
		.src_channel        (id_router_005_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                             //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_006 (
		.sink_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                      //       src.ready
		.src_valid          (id_router_006_src_valid),                                                      //          .valid
		.src_data           (id_router_006_src_data),                                                       //          .data
		.src_channel        (id_router_006_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                 //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_007 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                //          .valid
		.src_data           (id_router_007_src_data),                                                                 //          .data
		.src_channel        (id_router_007_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                           //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_008 (
		.sink_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                               //          .valid
		.src_data           (id_router_008_src_data),                                                //          .data
		.src_channel        (id_router_008_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                          //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_009 (
		.sink_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                      //          .valid
		.src_data           (id_router_009_src_data),                                                                       //          .data
		.src_channel        (id_router_009_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                                 //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_010 (
		.sink_ready         (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (remote_update_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                     //       src.ready
		.src_valid          (id_router_010_src_valid),                                                     //          .valid
		.src_data           (id_router_010_src_data),                                                      //          .data
		.src_channel        (id_router_010_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_011 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                     //       src.ready
		.src_valid          (id_router_011_src_valid),                                                     //          .valid
		.src_data           (id_router_011_src_data),                                                      //          .data
		.src_channel        (id_router_011_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_012 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                        //       src.ready
		.src_valid          (id_router_012_src_valid),                                                        //          .valid
		.src_data           (id_router_012_src_data),                                                         //          .data
		.src_channel        (id_router_012_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                   //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_005 id_router_013 (
		.sink_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                  //       src.ready
		.src_valid          (id_router_013_src_valid),                                                  //          .valid
		.src_data           (id_router_013_src_data),                                                   //          .data
		.src_channel        (id_router_013_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                             //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_addr_router_004 addr_router_004 (
		.sink_ready         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                                    // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                                             //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                                             //          .valid
		.src_data           (addr_router_004_src_data),                                                                              //          .data
		.src_channel        (addr_router_004_src_channel),                                                                           //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                                        //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_014 id_router_014 (
		.sink_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                  //       src.ready
		.src_valid          (id_router_014_src_valid),                                                  //          .valid
		.src_data           (id_router_014_src_data),                                                   //          .data
		.src_channel        (id_router_014_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                             //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_id_router_015 id_router_015 (
		.sink_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                           //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                              //       src.ready
		.src_valid          (id_router_015_src_valid),                                              //          .valid
		.src_data           (id_router_015_src_data),                                               //          .data
		.src_channel        (id_router_015_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                         //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (80),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (87),
		.PKT_TRANS_POSTED          (65),
		.PKT_TRANS_WRITE           (66),
		.MAX_OUTSTANDING_RESPONSES (72),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (70),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (70),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.MAX_OUTSTANDING_RESPONSES (6),
		.PIPELINED                 (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (pll_c2_out),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_003 (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_004_src_data),           //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_004_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_004_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_004_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_004_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (pll_c0_out),                          //       cr0.clk
		.reset                 (rst_controller_003_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),         //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),          //          .data
		.sink0_channel         (width_adapter_002_src_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                          // reset_in0.reset
		.reset_in1  (~ddr_sdram_reset_request_n_reset),  // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk),                               //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~ddr_sdram_reset_request_n_reset),   // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (pll_c2_out),                         //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~ddr_sdram_reset_request_n_reset),   // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (pll_c3_out),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~ddr_sdram_reset_request_n_reset),   // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (pll_c0_out),                         //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~ddr_sdram_reset_request_n_reset),   // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (ddr_sdram_phy_clk_out),              //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (clk),                                //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pll_c0_out),                         //        clk.clk
		.reset              (rst_controller_003_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)     //           .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //           .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pll_c0_out),                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (ddr_sdram_phy_clk_out),                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (ddr_sdram_phy_clk_out),                 //       clk.clk
		.reset              (~ddr_sdram_reset_request_n_reset),      // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (pll_c2_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_003_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_003_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_003_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_003_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_003_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_003_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_003_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_003_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_003_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_003_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_003_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_003_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_003_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_003_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_003_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_003_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_003_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_003_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_003_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_003_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_003_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_003_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_003_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_003_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_003_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_003_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_003_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_003_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_003_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_003_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_003_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_003_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_003_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_003_src7_endofpacket),   //           .endofpacket
		.src8_ready         (cmd_xbar_demux_003_src8_ready),         //       src8.ready
		.src8_valid         (cmd_xbar_demux_003_src8_valid),         //           .valid
		.src8_data          (cmd_xbar_demux_003_src8_data),          //           .data
		.src8_channel       (cmd_xbar_demux_003_src8_channel),       //           .channel
		.src8_startofpacket (cmd_xbar_demux_003_src8_startofpacket), //           .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_003_src8_endofpacket)    //           .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_006 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_007 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_008 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_009 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_010 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_011 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_012 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_005 rsp_xbar_demux_013 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_005_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_006_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_007_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_008_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_009_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (crosser_003_out_ready),                 //     sink5.ready
		.sink5_valid         (crosser_003_out_valid),                 //          .valid
		.sink5_channel       (crosser_003_out_channel),               //          .channel
		.sink5_data          (crosser_003_out_data),                  //          .data
		.sink5_startofpacket (crosser_003_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket   (crosser_003_out_endofpacket),           //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_011_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (crosser_004_out_ready),                 //     sink7.ready
		.sink7_valid         (crosser_004_out_valid),                 //          .valid
		.sink7_channel       (crosser_004_out_channel),               //          .channel
		.sink7_data          (crosser_004_out_data),                  //          .data
		.sink7_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink7_endofpacket   (crosser_004_out_endofpacket),           //          .endofpacket
		.sink8_ready         (crosser_005_out_ready),                 //     sink8.ready
		.sink8_valid         (crosser_005_out_valid),                 //          .valid
		.sink8_channel       (crosser_005_out_channel),               //          .channel
		.sink8_data          (crosser_005_out_data),                  //          .data
		.sink8_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink8_endofpacket   (crosser_005_out_endofpacket)            //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_003_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_003_cmd_src_channel),           //           .channel
		.sink_data          (limiter_003_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_003_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_003_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_003_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_004_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_004_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_004_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_004_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_004_src1_endofpacket)    //           .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_014 rsp_xbar_demux_014 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_demux_014 rsp_xbar_demux_015 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	cycloneIII_3c25_niosII_standard_sopc_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_014_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_015_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (74),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (77),
		.IN_PKT_BURST_SIZE_L           (75),
		.IN_PKT_RESPONSE_STATUS_H      (95),
		.IN_PKT_RESPONSE_STATUS_L      (94),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (79),
		.IN_PKT_BURST_TYPE_L           (78),
		.IN_ST_DATA_W                  (96),
		.OUT_PKT_ADDR_H                (96),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (106),
		.OUT_PKT_BYTE_CNT_L            (103),
		.OUT_PKT_TRANS_COMPRESSED_READ (97),
		.OUT_PKT_BURST_SIZE_H          (113),
		.OUT_PKT_BURST_SIZE_L          (111),
		.OUT_PKT_RESPONSE_STATUS_H     (131),
		.OUT_PKT_RESPONSE_STATUS_L     (130),
		.OUT_PKT_TRANS_EXCLUSIVE       (102),
		.OUT_PKT_BURST_TYPE_H          (115),
		.OUT_PKT_BURST_TYPE_L          (114),
		.OUT_ST_DATA_W                 (132),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (ddr_sdram_phy_clk_out),                 //       clk.clk
		.reset                (~ddr_sdram_reset_request_n_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data             (width_adapter_src_data),                //          .data
		.out_channel          (width_adapter_src_channel),             //          .channel
		.out_valid            (width_adapter_src_valid),               //          .valid
		.out_ready            (width_adapter_src_ready),               //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),       //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (96),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (106),
		.IN_PKT_BYTE_CNT_L             (103),
		.IN_PKT_TRANS_COMPRESSED_READ  (97),
		.IN_PKT_BURSTWRAP_H            (110),
		.IN_PKT_BURSTWRAP_L            (107),
		.IN_PKT_BURST_SIZE_H           (113),
		.IN_PKT_BURST_SIZE_L           (111),
		.IN_PKT_RESPONSE_STATUS_H      (131),
		.IN_PKT_RESPONSE_STATUS_L      (130),
		.IN_PKT_TRANS_EXCLUSIVE        (102),
		.IN_PKT_BURST_TYPE_H           (115),
		.IN_PKT_BURST_TYPE_L           (114),
		.IN_ST_DATA_W                  (132),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (77),
		.OUT_PKT_BURST_SIZE_L          (75),
		.OUT_PKT_RESPONSE_STATUS_H     (95),
		.OUT_PKT_RESPONSE_STATUS_L     (94),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (79),
		.OUT_PKT_BURST_TYPE_L          (78),
		.OUT_ST_DATA_W                 (96),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (ddr_sdram_phy_clk_out),               //       clk.clk
		.reset                (~ddr_sdram_reset_request_n_reset),    // clk_reset.reset
		.in_valid             (id_router_004_src_valid),             //      sink.valid
		.in_channel           (id_router_004_src_channel),           //          .channel
		.in_startofpacket     (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_004_src_ready),             //          .ready
		.in_data              (id_router_004_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (93),
		.IN_PKT_RESPONSE_STATUS_L      (92),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (94),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (75),
		.OUT_PKT_RESPONSE_STATUS_L     (74),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (76),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_004_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_004_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_004_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_004_src0_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (75),
		.IN_PKT_RESPONSE_STATUS_L      (74),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (76),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (93),
		.OUT_PKT_RESPONSE_STATUS_L     (92),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (94),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (pll_c0_out),                          //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_014_src_valid),             //      sink.valid
		.in_channel           (id_router_014_src_channel),           //          .channel
		.in_startofpacket     (id_router_014_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_014_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_014_src_ready),             //          .ready
		.in_data              (id_router_014_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c3_out),                            //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_003_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_003_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_003_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_003_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_003_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_003_src5_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c0_out),                            //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_003_src7_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_003_src7_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_003_src7_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_003_src7_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_003_src7_channel),       //              .channel
		.in_data           (cmd_xbar_demux_003_src7_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_005_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_003_src8_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_003_src8_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_003_src8_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_003_src8_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_003_src8_channel),       //              .channel
		.in_data           (cmd_xbar_demux_003_src8_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (pll_c3_out),                            //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_010_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_010_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_010_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_010_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (pll_c0_out),                            //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (9),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_005_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_013_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_013_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_013_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_013_src0_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	cycloneIII_3c25_niosII_standard_sopc_irq_mapper irq_mapper (
		.clk           (pll_c0_out),                         //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

endmodule
