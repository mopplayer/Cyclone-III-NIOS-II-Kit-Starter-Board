/* cycloneIII_3c25_start_golden_top.v
 This is a top level wrapper file that instanciates the
 golden top project

*/
module cycloneIII_3c25_start_golden_top(

// global signals:
input            osc_clk,
input            reset_n,

// the_button and led pios
input   [  3: 0] button,
output  [  3: 0] led, 		// note: led[1] needs distinct Assignment Setting: 
							// I/O Standard = "SSTL-2 Class I" 
							// due to location within the DDR block  
													              
// ddr
output  [ 12: 0] ddr_addr,
output  [  1: 0] ddr_ba,
output           ddr_cas_n,
output           ddr_cke,
inout            ddr_clk_n,
inout            ddr_clk,
output           ddr_cs_n,
output  [  1: 0] ddr_dm,
inout   [ 15: 0] ddr_dq,
inout   [  1: 0] ddr_dqs,
output           ddr_ras_n,
output           ddr_we_n,
                 
// flash/ssram shared bus
output  [ 23: 0] flash_ssram_a,
output			 flash_ssram_a24,		//to support 32MBytes & 64MBytes flash 
output			 flash_ssram_a25,		//to support 32MBytes & 64MBytes flash 
inout   [ 31: 0] flash_ssram_d,                             
               
output           ssram_adsc_n,
output  [  3: 0] ssram_bw_n,
output           ssram_bwe_n,
output           ssram_ce_n,
output           ssram_oe_n,
output           flash_oe_n,
output           flash_cs_n,
output           flash_wr_n,
output           ssram_clk,
output           flash_reset_n,           
                                  
//output           hsmc_clk,


// LCD Multimedia HSMC
inout	HC_ADC_BUSY,
output 			HC_ADC_CS_N,
output 			HC_ADC_DCLK,
output 			HC_ADC_DIN,
input			HC_ADC_DOUT,
input			HC_ADC_PENIRQ_N,
input		HC_AUD_ADCDAT,
inout		HC_AUD_ADCLRCK,
inout		HC_AUD_BCLK,
inout		HC_AUD_DACDAT,
inout		HC_AUD_DACLRCK,
inout		HC_AUD_XCK,
output			HC_DEN,
output			HC_ETH_RESET_N,
inout		HC_GREST,
output			HC_HD,
inout		HC_I2C_SCLK,
inout		HC_I2C_SDAT,
inout			HC_ID_I2CDAT,
output			HC_ID_I2CSCL,
output  [  7: 0] HC_LCD_DATA,
output			HC_MDC,
inout			HC_MDIO,
inout		HC_NCLK,
inout		HC_PS2_CLK,
inout		HC_PS2_DAT,
input			HC_RX_CLK,
input			HC_RX_COL,
input			HC_RX_CRS,
input  [  3: 0] HC_RX_D,
input			HC_RX_DV,
input			HC_RX_ERR,
output			HC_SCEN,
output			HC_SD_CLK,
output			HC_SD_CMD,
input			HC_SD_DAT,
output			HC_SD_DAT3,
inout			HC_SDA,
input		HC_TD_27MHZ,
inout		HC_TD_D0,
inout		HC_TD_D1,
inout		HC_TD_D2,
inout		HC_TD_D3,
inout		HC_TD_D4,
inout		HC_TD_D5,
inout		HC_TD_D6,
inout		HC_TD_D7,
inout		HC_TD_HS,
inout		HC_TD_RESET,
inout		HC_TD_VS,
input			HC_TX_CLK,
output [  3: 0] HC_TX_D,
output			HC_TX_EN,
inout		HC_UART_RXD,
inout		HC_UART_TXD,
output			HC_VD,
inout		HC_VGA_BLANK,
inout		HC_VGA_CLOCK,
inout  [   9:0]	HC_VGA_DATA,
inout		HC_VGA_HS,
inout		HC_VGA_SYNC,
inout		HC_VGA_VS

			
				
/* hsmc
input 	hsmc_clkin0,
input	hsmc_clkin_n1,
input	hsmc_clkin_n2,
input	hsmc_clkin_p1,
input 	hsmc_clkin_p2,
output  hsmc_clkout0,
output	hsmc_clkout_n1,
output	hsmc_clkout_n2,
output	hsmc_clkout_p1,
output	hsmc_clkout_p2,
inout 	hsmc_d0,
inout	hsmc_d1,
inout	hsmc_d2,
inout	hsmc_d3,
inout	hsmc_d4,
inout	hsmc_d5,
inout	hsmc_d6,
inout	hsmc_d7,
inout	hsmc_d8,
inout	hsmc_d9,
inout	hsmc_d10,
inout	hsmc_d11,
inout	hsmc_d12,
inout	hsmc_d13,
inout	hsmc_d14,
inout	hsmc_d15,
inout	hsmc_d16,
inout	hsmc_d17,
inout	hsmc_d18,
inout	hsmc_d19,
inout	hsmc_rx_n4,
inout	hsmc_rx_n5,
inout	hsmc_rx_n6,
inout	hsmc_rx_n7,
inout	hsmc_rx_n8,
inout	hsmc_rx_n9,
inout	hsmc_rx_n10,
inout	hsmc_rx_n11,
inout	hsmc_rx_n12,
inout	hsmc_rx_n13,
inout	hsmc_rx_n14,
inout	hsmc_rx_n15,
inout	hsmc_rx_n16,
inout	hsmc_rx_p4,
inout	hsmc_rx_p5,
inout	hsmc_rx_p6,
inout	hsmc_rx_p7,
inout	hsmc_rx_p8,
inout	hsmc_rx_p9,
inout	hsmc_rx_p10,
inout	hsmc_rx_p11,
inout	hsmc_rx_p12,
inout	hsmc_rx_p13,
inout	hsmc_rx_p14,
inout	hsmc_rx_p15,
inout	hsmc_rx_p16,
inout	hsmc_scl,
inout	hsmc_sda,
inout	hsmc_tx_n4,
inout	hsmc_tx_n5,
inout	hsmc_tx_n6,
inout	hsmc_tx_n7,
inout	hsmc_tx_n8,
inout	hsmc_tx_n9,
inout	hsmc_tx_n10,
inout	hsmc_tx_n11,
inout	hsmc_tx_n12,
inout	hsmc_tx_n13,
inout	hsmc_tx_n14,
inout	hsmc_tx_n15,
inout	hsmc_tx_n16,
inout	hsmc_tx_p4,
inout	hsmc_tx_p5,
inout	hsmc_tx_p6,
inout	hsmc_tx_p7,
inout	hsmc_tx_p8,
inout	hsmc_tx_p9,
inout	hsmc_tx_p10,
inout	hsmc_tx_p11,
inout	hsmc_tx_p12,
inout	hsmc_tx_p13,
inout	hsmc_tx_p14,
inout	hsmc_tx_p15,
inout	hsmc_tx_p16		*/
								
);  
endmodule
