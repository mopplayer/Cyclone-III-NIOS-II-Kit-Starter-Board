//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2012 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arbitrator (
                                                                                                  // inputs:
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n,
                                                                                                   clk,
                                                                                                   cpu_data_master_address_to_slave,
                                                                                                   cpu_data_master_latency_counter,
                                                                                                   cpu_data_master_read,
                                                                                                   cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
                                                                                                   cpu_data_master_write,
                                                                                                   cpu_data_master_writedata,
                                                                                                   reset_n,

                                                                                                  // outputs:
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write,
                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata,
                                                                                                   cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                                                                                   cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                                                                                   cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                                                                                   cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                                                                                   d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer
                                                                                                )
;

  output  [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa;
  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write;
  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata;
  output           cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  output           cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  output           cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  output           cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  output           d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n;
  input            clk;
  input   [ 27: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;

  wire    [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_allgrants;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_allow_new_arb_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_bursting_master_saved_grant;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_counter_enable;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter_next_value;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_set_values;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_beginbursttransfer_internal;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_begins_xfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_grant_vector;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_read_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_write_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_master_qreq_vector;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_non_bursting_master_requests;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reg_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_unreg_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_read;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_write;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata;
  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_saved_grant_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  reg              d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 27: 0] shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_from_cpu_data_master;
  wire             wait_for_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
    end


  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0));
  //assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata;

  assign cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 = ({cpu_data_master_address_to_slave[27 : 6] , 6'b0} == 28'h8000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter set values, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_set_values = 1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_non_bursting_master_requests mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_non_bursting_master_requests = cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_bursting_master_saved_grant mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_bursting_master_saved_grant = 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter_next_value assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter_next_value = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_firsttransfer ? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_set_values - 1) : |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter ? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter - 1) : 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_allgrants all slave grants, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_allgrants = |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_grant_vector;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer = ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_read | accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_write);

  //end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer & (~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter arbitration counter enable, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_counter_enable = (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_allgrants) | (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_non_bursting_master_requests);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter <= 0;
      else if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_counter_enable)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable <= 0;
      else if ((|accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_master_qreq_vector & end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0) | (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_non_bursting_master_requests))
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable <= |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter_next_value;
    end


  //cpu/data_master accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/cpu_interface0 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable & cpu_data_master_continuerequest;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable2 = |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arb_share_counter_next_value;

  //cpu/data_master accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/cpu_interface0 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_continuerequest at least one master continues requesting, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 = cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0, which is an e_mux
  assign cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 = cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & cpu_data_master_read & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_read;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 = cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;

  //cpu/data_master saved-grant accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/cpu_interface0, which is an e_assign
  assign cpu_data_master_saved_grant_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 = cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;

  //allow new arb cycle for accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/cpu_interface0, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_master_qreq_vector = 1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n = reset_n;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect = cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_firsttransfer first transaction, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_firsttransfer = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_begins_xfer ? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_unreg_firsttransfer : accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reg_firsttransfer;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_unreg_firsttransfer first transaction, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_unreg_firsttransfer = ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_any_continuerequest);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reg_firsttransfer <= 1'b1;
      else if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_begins_xfer)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reg_firsttransfer <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_unreg_firsttransfer;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_beginbursttransfer_internal = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_begins_xfer;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write assignment, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write = cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & cpu_data_master_write;

  assign shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_from_cpu_data_master = cpu_data_master_address_to_slave;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address = shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_from_cpu_data_master >> 2;

  //d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer <= 1;
      else 
        d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_read in a cycle, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_read = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_read_cycle & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_read_cycle assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_read_cycle = cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_read_cycle;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_write in a cycle, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waits_for_write = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_write_cycle & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_write_cycle assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_write_cycle = cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_in_a_write_cycle;

  assign wait_for_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_counter = 0;
  //assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/cpu_interface0 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arbitrator (
                                                                                               // inputs:
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata,
                                                                                                clk,
                                                                                                reset_n,

                                                                                               // outputs:
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect,
                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa,
                                                                                                d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer
                                                                                             )
;

  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect;
  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa;
  output           d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata;
  input            clk;
  input            reset_n;

  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_arbiterlock;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_arbiterlock2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_saved_grant_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_allgrants;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_allow_new_arb_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_bursting_master_saved_grant;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_counter_enable;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter_next_value;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_set_values;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_beginbursttransfer_internal;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_begins_xfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_grant_vector;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_read_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_write_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_master_qreq_vector;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_non_bursting_master_requests;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_reg_firsttransfer;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_unreg_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_read;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_write;
  reg              d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 31: 0] shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master;
  wire             wait_for_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
    end


  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_begins_xfer = ~d1_reasons_to_wait & ((accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave));
  //assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave = ({accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave[31 : 3] , 3'b0} == 32'h0) & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write);
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter set values, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_set_values = 1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_non_bursting_master_requests mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_non_bursting_master_requests = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_bursting_master_saved_grant = 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter_next_value = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_firsttransfer ? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_set_values - 1) : |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter ? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter - 1) : 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_allgrants all slave grants, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_allgrants = |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_grant_vector;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer = ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_read | accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer & (~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_allgrants) | (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_non_bursting_master_requests);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter <= 0;
      else if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_counter_enable)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable <= 0;
      else if ((|accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_master_qreq_vector & end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave) | (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_non_bursting_master_requests))
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable <= |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_master accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_slave arbiterlock, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_arbiterlock = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_continuerequest;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable2 = |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arb_share_counter_next_value;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_master accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_slave arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_arbiterlock2 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_continuerequest;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_continuerequest = 1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_continuerequest continued request, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_continuerequest = 1;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  //master is always granted when requested
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_master saved-grant accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_slave, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_saved_grant_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;

  //allow new arb cycle for accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_slave, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_master_qreq_vector = 1;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_firsttransfer first transaction, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_firsttransfer = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_begins_xfer ? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_unreg_firsttransfer : accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_reg_firsttransfer;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_unreg_firsttransfer = ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_any_continuerequest);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_reg_firsttransfer <= 1'b1;
      else if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_begins_xfer)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_reg_firsttransfer <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_unreg_firsttransfer;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_beginbursttransfer_internal = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_begins_xfer;

  assign shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address = shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master >> 2;

  //d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer <= 1;
      else 
        d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_read in a cycle, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_read = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_read_cycle & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_begins_xfer;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_read_cycle assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_read_cycle = 0;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_read_cycle;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_write in a cycle, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_waits_for_write = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_write_cycle & 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_write_cycle assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_write_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_in_a_write_cycle;

  assign wait_for_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arbitrator (
                                                                                                               // inputs:
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n,
                                                                                                                clk,
                                                                                                                reset_n,

                                                                                                               // outputs:
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n,
                                                                                                                accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa,
                                                                                                                d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer
                                                                                                             )
;

  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read;
  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa;
  output           d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n;
  input            clk;
  input            reset_n;

  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_arbiterlock;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_arbiterlock2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_saved_grant_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_allgrants;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_allow_new_arb_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_bursting_master_saved_grant;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_counter_enable;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter_next_value;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_set_values;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_beginbursttransfer_internal;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begins_xfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_grant_vector;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_read_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_write_cycle;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_master_qreq_vector;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_non_bursting_master_requests;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reg_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_unreg_firsttransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_read;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_write;
  reg              d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 31: 0] shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0;
  wire             wait_for_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
    end


  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begins_xfer = ~d1_reasons_to_wait & ((accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0));
  //assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 = (({accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave[31 : 2] , 2'b0} == 32'h0) & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read)) & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;
  //assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter set values, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_set_values = 1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_non_bursting_master_requests mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_non_bursting_master_requests = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_bursting_master_saved_grant mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_bursting_master_saved_grant = 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter_next_value assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter_next_value = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_firsttransfer ? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_set_values - 1) : |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter ? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter - 1) : 0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_allgrants all slave grants, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_allgrants = |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_grant_vector;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer = ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_read | accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_write);

  //end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer & (~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter arbitration counter enable, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_counter_enable = (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_allgrants) | (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_non_bursting_master_requests);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter <= 0;
      else if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_counter_enable)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable <= 0;
      else if ((|accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_master_qreq_vector & end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0) | (end_xfer_arb_share_counter_term_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_non_bursting_master_requests))
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable <= |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/internal_master0 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/sub_hw_draw_int_mandelbrot0 arbiterlock, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_arbiterlock = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_continuerequest;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable2 = |accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arb_share_counter_next_value;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/internal_master0 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/sub_hw_draw_int_mandelbrot0 arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_arbiterlock2 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_continuerequest;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_continuerequest at least one master continues requesting, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_continuerequest = 1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_continuerequest continued request, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_continuerequest = 1;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  //master is always granted when requested
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/internal_master0 saved-grant accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/sub_hw_draw_int_mandelbrot0, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_saved_grant_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;

  //allow new arb cycle for accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/sub_hw_draw_int_mandelbrot0, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_master_qreq_vector = 1;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begins_xfer;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n = reset_n;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_firsttransfer first transaction, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_firsttransfer = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begins_xfer ? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_unreg_firsttransfer : accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reg_firsttransfer;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_unreg_firsttransfer first transaction, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_unreg_firsttransfer = ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_any_continuerequest);

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reg_firsttransfer <= 1'b1;
      else if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begins_xfer)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reg_firsttransfer <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_unreg_firsttransfer;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_beginbursttransfer_internal = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begins_xfer;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read assignment, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;

  assign shifted_address_to_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave;
  //d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer <= 1;
      else 
        d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_read in a cycle, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_read = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_read_cycle & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_read_cycle assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_read_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_read_cycle;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_write in a cycle, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waits_for_write = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_write_cycle & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_write_cycle assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_in_a_write_cycle;

  assign wait_for_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/sub_hw_draw_int_mandelbrot0 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbitrator (
                                                                                                                                                  // inputs:
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2,
                                                                                                                                                   clk,
                                                                                                                                                   colour_lookup_table_s2_readdata_from_sa,
                                                                                                                                                   d1_colour_lookup_table_s2_end_xfer,
                                                                                                                                                   reset_n,

                                                                                                                                                  // outputs:
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n
                                                                                                                                                )
;

  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter;
  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2;
  input            clk;
  input   [ 31: 0] colour_lookup_table_s2_readdata_from_sa;
  input            d1_colour_lookup_table_s2_end_xfer;
  input            reset_n;

  reg     [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_last_time;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_is_granted_some_slave;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_but_no_slave_selected;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_last_time;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run_delayed;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n;
  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter;
  wire             pre_flush_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2 | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2) & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2 | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2) & ((~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2 | ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read) | (1 & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read))));

  //cascaded wait assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave = {22'b10001000000000111,
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address[9 : 0]};

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_but_no_slave_selected <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_but_no_slave_selected <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_is_granted_some_slave = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2;

  //run delay, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run_delayed <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run_delayed <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run;
    end


  //The Flushificator, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush && accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run_delayed;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_but_no_slave_selected |
    (pre_flush_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid & ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified);

  //The Exported Flushificator, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 readdata mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata = colour_lookup_table_s2_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter <= p1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter = ((accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_run & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read))? latency_load_value :
    (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter)? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read);
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbitrator (
                                                                                                                                                  // inputs:
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata,
                                                                                                                                                   clk,
                                                                                                                                                   d1_frame_buffer_pipeline_bridge_s1_end_xfer,
                                                                                                                                                   frame_buffer_pipeline_bridge_s1_waitrequest_from_sa,
                                                                                                                                                   reset_n,

                                                                                                                                                  // outputs:
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave,
                                                                                                                                                   accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n
                                                                                                                                                )
;

  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address;
  input   [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata;
  input            clk;
  input            d1_frame_buffer_pipeline_bridge_s1_end_xfer;
  input            frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;
  input            reset_n;

  reg     [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_last_time;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave;
  reg     [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable_last_time;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_run;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write_last_time;
  reg     [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1 | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1) & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1 | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1) & ((~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1 | ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write) | (1 & ~frame_buffer_pipeline_bridge_s1_waitrequest_from_sa & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write))));

  //cascaded wait assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave = {7'b0,
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address[24 : 0]};

  //actual waitrequest port, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write);
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata_last_time) & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write)
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_arbitrator (
                                                                                                // inputs:
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address,
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave,
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave,
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave,
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write,
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata,
                                                                                                 clk,
                                                                                                 d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer,
                                                                                                 reset_n,

                                                                                                // outputs:
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave,
                                                                                                 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest
                                                                                              )
;

  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata;
  input            clk;
  input            d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
  input            reset_n;

  reg     [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_last_time;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_run;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write_last_time;
  reg     [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata_last_time;
  reg              active_and_waiting_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & ((~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write | (1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write)));

  //cascaded wait assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave = {29'b0,
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address[2 : 0]};

  //actual waitrequest port, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest = ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/dummy_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write);
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata_last_time) & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write)
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_arbitrator (
                                                                                                    // inputs:
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa,
                                                                                                     clk,
                                                                                                     d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer,
                                                                                                     reset_n,

                                                                                                    // outputs:
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata,
                                                                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n
                                                                                                  )
;

  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave;
  output  [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa;
  input            clk;
  input            d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
  input            reset_n;

  reg     [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_last_time;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_last_time;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_run;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n;
  reg              active_and_waiting_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & ((~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 | ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read) | (1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read))));

  //cascaded wait assignment, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave = {30'b0,
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address[1 : 0]};

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/internal_master0 readdata mux, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/internal_master0 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read);
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_last_time <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_last_time <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read != accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_last_time))
        begin
          $write("%0d ns: accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_pipeline_bridge_m1_to_clock_crossing_bridge_s1_module (
                                                                            // inputs:
                                                                             clear_fifo,
                                                                             clk,
                                                                             data_in,
                                                                             read,
                                                                             reset_n,
                                                                             sync_reset,
                                                                             write,

                                                                            // outputs:
                                                                             data_out,
                                                                             empty,
                                                                             fifo_contains_ones_n,
                                                                             full
                                                                          )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  wire             full_16;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_15;
  assign empty = !full_0;
  assign full_16 = 0;
  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    0;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_bridge_s1_arbitrator (
                                             // inputs:
                                              clk,
                                              clock_crossing_bridge_s1_endofpacket,
                                              clock_crossing_bridge_s1_readdata,
                                              clock_crossing_bridge_s1_readdatavalid,
                                              clock_crossing_bridge_s1_waitrequest,
                                              pipeline_bridge_m1_address_to_slave,
                                              pipeline_bridge_m1_burstcount,
                                              pipeline_bridge_m1_byteenable,
                                              pipeline_bridge_m1_chipselect,
                                              pipeline_bridge_m1_latency_counter,
                                              pipeline_bridge_m1_read,
                                              pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                              pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                              pipeline_bridge_m1_write,
                                              pipeline_bridge_m1_writedata,
                                              reset_n,

                                             // outputs:
                                              clock_crossing_bridge_s1_address,
                                              clock_crossing_bridge_s1_byteenable,
                                              clock_crossing_bridge_s1_endofpacket_from_sa,
                                              clock_crossing_bridge_s1_nativeaddress,
                                              clock_crossing_bridge_s1_read,
                                              clock_crossing_bridge_s1_readdata_from_sa,
                                              clock_crossing_bridge_s1_reset_n,
                                              clock_crossing_bridge_s1_waitrequest_from_sa,
                                              clock_crossing_bridge_s1_write,
                                              clock_crossing_bridge_s1_writedata,
                                              d1_clock_crossing_bridge_s1_end_xfer,
                                              pipeline_bridge_m1_granted_clock_crossing_bridge_s1,
                                              pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1,
                                              pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1,
                                              pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                              pipeline_bridge_m1_requests_clock_crossing_bridge_s1
                                           )
;

  output  [  8: 0] clock_crossing_bridge_s1_address;
  output  [  3: 0] clock_crossing_bridge_s1_byteenable;
  output           clock_crossing_bridge_s1_endofpacket_from_sa;
  output  [  8: 0] clock_crossing_bridge_s1_nativeaddress;
  output           clock_crossing_bridge_s1_read;
  output  [ 31: 0] clock_crossing_bridge_s1_readdata_from_sa;
  output           clock_crossing_bridge_s1_reset_n;
  output           clock_crossing_bridge_s1_waitrequest_from_sa;
  output           clock_crossing_bridge_s1_write;
  output  [ 31: 0] clock_crossing_bridge_s1_writedata;
  output           d1_clock_crossing_bridge_s1_end_xfer;
  output           pipeline_bridge_m1_granted_clock_crossing_bridge_s1;
  output           pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1;
  output           pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1;
  output           pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  output           pipeline_bridge_m1_requests_clock_crossing_bridge_s1;
  input            clk;
  input            clock_crossing_bridge_s1_endofpacket;
  input   [ 31: 0] clock_crossing_bridge_s1_readdata;
  input            clock_crossing_bridge_s1_readdatavalid;
  input            clock_crossing_bridge_s1_waitrequest;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  wire    [  8: 0] clock_crossing_bridge_s1_address;
  wire             clock_crossing_bridge_s1_allgrants;
  wire             clock_crossing_bridge_s1_allow_new_arb_cycle;
  wire             clock_crossing_bridge_s1_any_bursting_master_saved_grant;
  wire             clock_crossing_bridge_s1_any_continuerequest;
  wire             clock_crossing_bridge_s1_arb_counter_enable;
  reg              clock_crossing_bridge_s1_arb_share_counter;
  wire             clock_crossing_bridge_s1_arb_share_counter_next_value;
  wire             clock_crossing_bridge_s1_arb_share_set_values;
  wire             clock_crossing_bridge_s1_beginbursttransfer_internal;
  wire             clock_crossing_bridge_s1_begins_xfer;
  wire    [  3: 0] clock_crossing_bridge_s1_byteenable;
  wire             clock_crossing_bridge_s1_end_xfer;
  wire             clock_crossing_bridge_s1_endofpacket_from_sa;
  wire             clock_crossing_bridge_s1_firsttransfer;
  wire             clock_crossing_bridge_s1_grant_vector;
  wire             clock_crossing_bridge_s1_in_a_read_cycle;
  wire             clock_crossing_bridge_s1_in_a_write_cycle;
  wire             clock_crossing_bridge_s1_master_qreq_vector;
  wire             clock_crossing_bridge_s1_move_on_to_next_transaction;
  wire    [  8: 0] clock_crossing_bridge_s1_nativeaddress;
  wire             clock_crossing_bridge_s1_non_bursting_master_requests;
  wire             clock_crossing_bridge_s1_read;
  wire    [ 31: 0] clock_crossing_bridge_s1_readdata_from_sa;
  wire             clock_crossing_bridge_s1_readdatavalid_from_sa;
  reg              clock_crossing_bridge_s1_reg_firsttransfer;
  wire             clock_crossing_bridge_s1_reset_n;
  reg              clock_crossing_bridge_s1_slavearbiterlockenable;
  wire             clock_crossing_bridge_s1_slavearbiterlockenable2;
  wire             clock_crossing_bridge_s1_unreg_firsttransfer;
  wire             clock_crossing_bridge_s1_waitrequest_from_sa;
  wire             clock_crossing_bridge_s1_waits_for_read;
  wire             clock_crossing_bridge_s1_waits_for_write;
  wire             clock_crossing_bridge_s1_write;
  wire    [ 31: 0] clock_crossing_bridge_s1_writedata;
  reg              d1_clock_crossing_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_clock_crossing_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_rdv_fifo_empty_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_rdv_fifo_output_from_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  wire             pipeline_bridge_m1_requests_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_saved_grant_clock_crossing_bridge_s1;
  wire    [ 26: 0] shifted_address_to_clock_crossing_bridge_s1_from_pipeline_bridge_m1;
  wire             wait_for_clock_crossing_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~clock_crossing_bridge_s1_end_xfer;
    end


  assign clock_crossing_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1));
  //assign clock_crossing_bridge_s1_readdata_from_sa = clock_crossing_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_bridge_s1_readdata_from_sa = clock_crossing_bridge_s1_readdata;

  assign pipeline_bridge_m1_requests_clock_crossing_bridge_s1 = ({pipeline_bridge_m1_address_to_slave[26 : 11] , 11'b0} == 27'h4000000) & pipeline_bridge_m1_chipselect;
  //assign clock_crossing_bridge_s1_waitrequest_from_sa = clock_crossing_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_bridge_s1_waitrequest_from_sa = clock_crossing_bridge_s1_waitrequest;

  //assign clock_crossing_bridge_s1_readdatavalid_from_sa = clock_crossing_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_bridge_s1_readdatavalid_from_sa = clock_crossing_bridge_s1_readdatavalid;

  //clock_crossing_bridge_s1_arb_share_counter set values, which is an e_mux
  assign clock_crossing_bridge_s1_arb_share_set_values = 1;

  //clock_crossing_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign clock_crossing_bridge_s1_non_bursting_master_requests = pipeline_bridge_m1_requests_clock_crossing_bridge_s1;

  //clock_crossing_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign clock_crossing_bridge_s1_any_bursting_master_saved_grant = 0;

  //clock_crossing_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign clock_crossing_bridge_s1_arb_share_counter_next_value = clock_crossing_bridge_s1_firsttransfer ? (clock_crossing_bridge_s1_arb_share_set_values - 1) : |clock_crossing_bridge_s1_arb_share_counter ? (clock_crossing_bridge_s1_arb_share_counter - 1) : 0;

  //clock_crossing_bridge_s1_allgrants all slave grants, which is an e_mux
  assign clock_crossing_bridge_s1_allgrants = |clock_crossing_bridge_s1_grant_vector;

  //clock_crossing_bridge_s1_end_xfer assignment, which is an e_assign
  assign clock_crossing_bridge_s1_end_xfer = ~(clock_crossing_bridge_s1_waits_for_read | clock_crossing_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_clock_crossing_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_clock_crossing_bridge_s1 = clock_crossing_bridge_s1_end_xfer & (~clock_crossing_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //clock_crossing_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign clock_crossing_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_clock_crossing_bridge_s1 & clock_crossing_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_clock_crossing_bridge_s1 & ~clock_crossing_bridge_s1_non_bursting_master_requests);

  //clock_crossing_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_s1_arb_share_counter <= 0;
      else if (clock_crossing_bridge_s1_arb_counter_enable)
          clock_crossing_bridge_s1_arb_share_counter <= clock_crossing_bridge_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|clock_crossing_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_clock_crossing_bridge_s1) | (end_xfer_arb_share_counter_term_clock_crossing_bridge_s1 & ~clock_crossing_bridge_s1_non_bursting_master_requests))
          clock_crossing_bridge_s1_slavearbiterlockenable <= |clock_crossing_bridge_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 clock_crossing_bridge/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = clock_crossing_bridge_s1_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //clock_crossing_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_s1_slavearbiterlockenable2 = |clock_crossing_bridge_s1_arb_share_counter_next_value;

  //pipeline_bridge/m1 clock_crossing_bridge/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = clock_crossing_bridge_s1_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //clock_crossing_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign clock_crossing_bridge_s1_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1 = pipeline_bridge_m1_requests_clock_crossing_bridge_s1 & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0) | (1 < pipeline_bridge_m1_latency_counter) | (|pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register))));
  //unique name for clock_crossing_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign clock_crossing_bridge_s1_move_on_to_next_transaction = clock_crossing_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_pipeline_bridge_m1_to_clock_crossing_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pipeline_bridge_m1_to_clock_crossing_bridge_s1_module rdv_fifo_for_pipeline_bridge_m1_to_clock_crossing_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pipeline_bridge_m1_granted_clock_crossing_bridge_s1),
      .data_out             (pipeline_bridge_m1_rdv_fifo_output_from_clock_crossing_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (pipeline_bridge_m1_rdv_fifo_empty_clock_crossing_bridge_s1),
      .full                 (),
      .read                 (clock_crossing_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~clock_crossing_bridge_s1_waits_for_read)
    );

  assign pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register = ~pipeline_bridge_m1_rdv_fifo_empty_clock_crossing_bridge_s1;
  //local readdatavalid pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1 = clock_crossing_bridge_s1_readdatavalid_from_sa;

  //clock_crossing_bridge_s1_writedata mux, which is an e_mux
  assign clock_crossing_bridge_s1_writedata = pipeline_bridge_m1_writedata;

  //assign clock_crossing_bridge_s1_endofpacket_from_sa = clock_crossing_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clock_crossing_bridge_s1_endofpacket_from_sa = clock_crossing_bridge_s1_endofpacket;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_clock_crossing_bridge_s1 = pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1;

  //pipeline_bridge/m1 saved-grant clock_crossing_bridge/s1, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_clock_crossing_bridge_s1 = pipeline_bridge_m1_requests_clock_crossing_bridge_s1;

  //allow new arb cycle for clock_crossing_bridge/s1, which is an e_assign
  assign clock_crossing_bridge_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign clock_crossing_bridge_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign clock_crossing_bridge_s1_master_qreq_vector = 1;

  //clock_crossing_bridge_s1_reset_n assignment, which is an e_assign
  assign clock_crossing_bridge_s1_reset_n = reset_n;

  //clock_crossing_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_bridge_s1_firsttransfer = clock_crossing_bridge_s1_begins_xfer ? clock_crossing_bridge_s1_unreg_firsttransfer : clock_crossing_bridge_s1_reg_firsttransfer;

  //clock_crossing_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign clock_crossing_bridge_s1_unreg_firsttransfer = ~(clock_crossing_bridge_s1_slavearbiterlockenable & clock_crossing_bridge_s1_any_continuerequest);

  //clock_crossing_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (clock_crossing_bridge_s1_begins_xfer)
          clock_crossing_bridge_s1_reg_firsttransfer <= clock_crossing_bridge_s1_unreg_firsttransfer;
    end


  //clock_crossing_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign clock_crossing_bridge_s1_beginbursttransfer_internal = clock_crossing_bridge_s1_begins_xfer;

  //clock_crossing_bridge_s1_read assignment, which is an e_mux
  assign clock_crossing_bridge_s1_read = pipeline_bridge_m1_granted_clock_crossing_bridge_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //clock_crossing_bridge_s1_write assignment, which is an e_mux
  assign clock_crossing_bridge_s1_write = pipeline_bridge_m1_granted_clock_crossing_bridge_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_clock_crossing_bridge_s1_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //clock_crossing_bridge_s1_address mux, which is an e_mux
  assign clock_crossing_bridge_s1_address = shifted_address_to_clock_crossing_bridge_s1_from_pipeline_bridge_m1 >> 2;

  //slaveid clock_crossing_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign clock_crossing_bridge_s1_nativeaddress = pipeline_bridge_m1_address_to_slave >> 2;

  //d1_clock_crossing_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_clock_crossing_bridge_s1_end_xfer <= 1;
      else 
        d1_clock_crossing_bridge_s1_end_xfer <= clock_crossing_bridge_s1_end_xfer;
    end


  //clock_crossing_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign clock_crossing_bridge_s1_waits_for_read = clock_crossing_bridge_s1_in_a_read_cycle & clock_crossing_bridge_s1_waitrequest_from_sa;

  //clock_crossing_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign clock_crossing_bridge_s1_in_a_read_cycle = pipeline_bridge_m1_granted_clock_crossing_bridge_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = clock_crossing_bridge_s1_in_a_read_cycle;

  //clock_crossing_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign clock_crossing_bridge_s1_waits_for_write = clock_crossing_bridge_s1_in_a_write_cycle & clock_crossing_bridge_s1_waitrequest_from_sa;

  //clock_crossing_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign clock_crossing_bridge_s1_in_a_write_cycle = pipeline_bridge_m1_granted_clock_crossing_bridge_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = clock_crossing_bridge_s1_in_a_write_cycle;

  assign wait_for_clock_crossing_bridge_s1_counter = 0;
  //clock_crossing_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign clock_crossing_bridge_s1_byteenable = (pipeline_bridge_m1_granted_clock_crossing_bridge_s1)? pipeline_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_clock_crossing_bridge_s1 && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave clock_crossing_bridge/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_bridge_m1_arbitrator (
                                             // inputs:
                                              clk,
                                              clock_crossing_bridge_m1_address,
                                              clock_crossing_bridge_m1_byteenable,
                                              clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
                                              clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1,
                                              clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1,
                                              clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1,
                                              clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1,
                                              clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1,
                                              clock_crossing_bridge_m1_granted_push_buttons_s1,
                                              clock_crossing_bridge_m1_granted_sysid_control_slave,
                                              clock_crossing_bridge_m1_granted_system_tick_s1,
                                              clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1,
                                              clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port,
                                              clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                              clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1,
                                              clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1,
                                              clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1,
                                              clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1,
                                              clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1,
                                              clock_crossing_bridge_m1_qualified_request_push_buttons_s1,
                                              clock_crossing_bridge_m1_qualified_request_sysid_control_slave,
                                              clock_crossing_bridge_m1_qualified_request_system_tick_s1,
                                              clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1,
                                              clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port,
                                              clock_crossing_bridge_m1_read,
                                              clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                              clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1,
                                              clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1,
                                              clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1,
                                              clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1,
                                              clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1,
                                              clock_crossing_bridge_m1_read_data_valid_push_buttons_s1,
                                              clock_crossing_bridge_m1_read_data_valid_sysid_control_slave,
                                              clock_crossing_bridge_m1_read_data_valid_system_tick_s1,
                                              clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1,
                                              clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port,
                                              clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
                                              clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1,
                                              clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1,
                                              clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1,
                                              clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1,
                                              clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1,
                                              clock_crossing_bridge_m1_requests_push_buttons_s1,
                                              clock_crossing_bridge_m1_requests_sysid_control_slave,
                                              clock_crossing_bridge_m1_requests_system_tick_s1,
                                              clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1,
                                              clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port,
                                              clock_crossing_bridge_m1_write,
                                              clock_crossing_bridge_m1_writedata,
                                              d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                              d1_lcd_i2c_cs_s1_end_xfer,
                                              d1_lcd_i2c_dat_s1_end_xfer,
                                              d1_lcd_i2c_scl_s1_end_xfer,
                                              d1_pio_id_eeprom_dat_s1_end_xfer,
                                              d1_pio_id_eeprom_scl_s1_end_xfer,
                                              d1_push_buttons_s1_end_xfer,
                                              d1_sysid_control_slave_end_xfer,
                                              d1_system_tick_s1_end_xfer,
                                              d1_touchPanel_irq_n_s1_end_xfer,
                                              d1_touchPanel_spi_spi_control_port_end_xfer,
                                              jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                              jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                              lcd_i2c_cs_s1_readdata_from_sa,
                                              lcd_i2c_dat_s1_readdata_from_sa,
                                              lcd_i2c_scl_s1_readdata_from_sa,
                                              pio_id_eeprom_dat_s1_readdata_from_sa,
                                              pio_id_eeprom_scl_s1_readdata_from_sa,
                                              push_buttons_s1_readdata_from_sa,
                                              reset_n,
                                              sysid_control_slave_readdata_from_sa,
                                              system_tick_s1_readdata_from_sa,
                                              touchPanel_irq_n_s1_readdata_from_sa,
                                              touchPanel_spi_spi_control_port_endofpacket_from_sa,
                                              touchPanel_spi_spi_control_port_readdata_from_sa,

                                             // outputs:
                                              clock_crossing_bridge_m1_address_to_slave,
                                              clock_crossing_bridge_m1_endofpacket,
                                              clock_crossing_bridge_m1_latency_counter,
                                              clock_crossing_bridge_m1_readdata,
                                              clock_crossing_bridge_m1_readdatavalid,
                                              clock_crossing_bridge_m1_reset_n,
                                              clock_crossing_bridge_m1_waitrequest
                                           )
;

  output  [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  output           clock_crossing_bridge_m1_endofpacket;
  output           clock_crossing_bridge_m1_latency_counter;
  output  [ 31: 0] clock_crossing_bridge_m1_readdata;
  output           clock_crossing_bridge_m1_readdatavalid;
  output           clock_crossing_bridge_m1_reset_n;
  output           clock_crossing_bridge_m1_waitrequest;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address;
  input   [  3: 0] clock_crossing_bridge_m1_byteenable;
  input            clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  input            clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1;
  input            clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1;
  input            clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1;
  input            clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1;
  input            clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1;
  input            clock_crossing_bridge_m1_granted_push_buttons_s1;
  input            clock_crossing_bridge_m1_granted_sysid_control_slave;
  input            clock_crossing_bridge_m1_granted_system_tick_s1;
  input            clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1;
  input            clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port;
  input            clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  input            clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1;
  input            clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1;
  input            clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1;
  input            clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1;
  input            clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1;
  input            clock_crossing_bridge_m1_qualified_request_push_buttons_s1;
  input            clock_crossing_bridge_m1_qualified_request_sysid_control_slave;
  input            clock_crossing_bridge_m1_qualified_request_system_tick_s1;
  input            clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1;
  input            clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1;
  input            clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1;
  input            clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1;
  input            clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1;
  input            clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1;
  input            clock_crossing_bridge_m1_read_data_valid_push_buttons_s1;
  input            clock_crossing_bridge_m1_read_data_valid_sysid_control_slave;
  input            clock_crossing_bridge_m1_read_data_valid_system_tick_s1;
  input            clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1;
  input            clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port;
  input            clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  input            clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1;
  input            clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1;
  input            clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1;
  input            clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1;
  input            clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1;
  input            clock_crossing_bridge_m1_requests_push_buttons_s1;
  input            clock_crossing_bridge_m1_requests_sysid_control_slave;
  input            clock_crossing_bridge_m1_requests_system_tick_s1;
  input            clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1;
  input            clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input            d1_lcd_i2c_cs_s1_end_xfer;
  input            d1_lcd_i2c_dat_s1_end_xfer;
  input            d1_lcd_i2c_scl_s1_end_xfer;
  input            d1_pio_id_eeprom_dat_s1_end_xfer;
  input            d1_pio_id_eeprom_scl_s1_end_xfer;
  input            d1_push_buttons_s1_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_system_tick_s1_end_xfer;
  input            d1_touchPanel_irq_n_s1_end_xfer;
  input            d1_touchPanel_spi_spi_control_port_end_xfer;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] lcd_i2c_cs_s1_readdata_from_sa;
  input   [ 31: 0] lcd_i2c_dat_s1_readdata_from_sa;
  input   [ 31: 0] lcd_i2c_scl_s1_readdata_from_sa;
  input   [ 31: 0] pio_id_eeprom_dat_s1_readdata_from_sa;
  input   [ 31: 0] pio_id_eeprom_scl_s1_readdata_from_sa;
  input   [ 31: 0] push_buttons_s1_readdata_from_sa;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 15: 0] system_tick_s1_readdata_from_sa;
  input   [ 31: 0] touchPanel_irq_n_s1_readdata_from_sa;
  input            touchPanel_spi_spi_control_port_endofpacket_from_sa;
  input   [ 15: 0] touchPanel_spi_spi_control_port_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 10: 0] clock_crossing_bridge_m1_address_last_time;
  wire    [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  reg     [  3: 0] clock_crossing_bridge_m1_byteenable_last_time;
  wire             clock_crossing_bridge_m1_endofpacket;
  wire             clock_crossing_bridge_m1_is_granted_some_slave;
  reg              clock_crossing_bridge_m1_latency_counter;
  reg              clock_crossing_bridge_m1_read_but_no_slave_selected;
  reg              clock_crossing_bridge_m1_read_last_time;
  wire    [ 31: 0] clock_crossing_bridge_m1_readdata;
  wire             clock_crossing_bridge_m1_readdatavalid;
  wire             clock_crossing_bridge_m1_reset_n;
  wire             clock_crossing_bridge_m1_run;
  wire             clock_crossing_bridge_m1_waitrequest;
  reg              clock_crossing_bridge_m1_write_last_time;
  reg     [ 31: 0] clock_crossing_bridge_m1_writedata_last_time;
  wire             latency_load_value;
  wire             p1_clock_crossing_bridge_m1_latency_counter;
  wire             pre_flush_clock_crossing_bridge_m1_readdatavalid;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave) & ((~clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~(clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write)))) & ((~clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~(clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write)))) & 1 & (clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1 | ~clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1) & ((~clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_lcd_i2c_cs_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1 | ~clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1) & ((~clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_lcd_i2c_dat_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1 | ~clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1) & ((~clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_lcd_i2c_scl_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1 | ~clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1) & ((~clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_pio_id_eeprom_dat_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write)));

  //cascaded wait assignment, which is an e_assign
  assign clock_crossing_bridge_m1_run = r_1 & r_2 & r_3;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1 | ~clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1) & ((~clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_pio_id_eeprom_scl_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_push_buttons_s1 | ~clock_crossing_bridge_m1_requests_push_buttons_s1) & ((~clock_crossing_bridge_m1_qualified_request_push_buttons_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_push_buttons_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_push_buttons_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_sysid_control_slave | ~clock_crossing_bridge_m1_requests_sysid_control_slave) & ((~clock_crossing_bridge_m1_qualified_request_sysid_control_slave | ~clock_crossing_bridge_m1_read | (1 & ~d1_sysid_control_slave_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_sysid_control_slave | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_system_tick_s1 | ~clock_crossing_bridge_m1_requests_system_tick_s1) & ((~clock_crossing_bridge_m1_qualified_request_system_tick_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_system_tick_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_system_tick_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write))) & 1 & (clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1 | ~clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1) & ((~clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1 | ~clock_crossing_bridge_m1_read | (1 & ~d1_touchPanel_irq_n_s1_end_xfer & clock_crossing_bridge_m1_read))) & ((~clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1 | ~clock_crossing_bridge_m1_write | (1 & clock_crossing_bridge_m1_write)));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port | ~clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port) & ((~clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port | ~(clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write) | (1 & ~d1_touchPanel_spi_spi_control_port_end_xfer & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write)))) & ((~clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port | ~(clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write) | (1 & ~d1_touchPanel_spi_spi_control_port_end_xfer & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign clock_crossing_bridge_m1_address_to_slave = {clock_crossing_bridge_m1_address[10 : 6],
    1'b0,
    clock_crossing_bridge_m1_address[4 : 0]};

  //clock_crossing_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_read_but_no_slave_selected <= 0;
      else 
        clock_crossing_bridge_m1_read_but_no_slave_selected <= clock_crossing_bridge_m1_read & clock_crossing_bridge_m1_run & ~clock_crossing_bridge_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign clock_crossing_bridge_m1_is_granted_some_slave = clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave |
    clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1 |
    clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1 |
    clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1 |
    clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1 |
    clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1 |
    clock_crossing_bridge_m1_granted_push_buttons_s1 |
    clock_crossing_bridge_m1_granted_sysid_control_slave |
    clock_crossing_bridge_m1_granted_system_tick_s1 |
    clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1 |
    clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_clock_crossing_bridge_m1_readdatavalid = 0;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign clock_crossing_bridge_m1_readdatavalid = clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_push_buttons_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_sysid_control_slave |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_system_tick_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1 |
    clock_crossing_bridge_m1_read_but_no_slave_selected |
    pre_flush_clock_crossing_bridge_m1_readdatavalid |
    clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port;

  //clock_crossing_bridge/m1 readdata mux, which is an e_mux
  assign clock_crossing_bridge_m1_readdata = ({32 {~(clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave & clock_crossing_bridge_m1_read)}} | jtag_uart_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1 & clock_crossing_bridge_m1_read)}} | lcd_i2c_cs_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1 & clock_crossing_bridge_m1_read)}} | lcd_i2c_dat_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1 & clock_crossing_bridge_m1_read)}} | lcd_i2c_scl_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1 & clock_crossing_bridge_m1_read)}} | pio_id_eeprom_dat_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1 & clock_crossing_bridge_m1_read)}} | pio_id_eeprom_scl_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_push_buttons_s1 & clock_crossing_bridge_m1_read)}} | push_buttons_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_sysid_control_slave & clock_crossing_bridge_m1_read)}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_system_tick_s1 & clock_crossing_bridge_m1_read)}} | system_tick_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1 & clock_crossing_bridge_m1_read)}} | touchPanel_irq_n_s1_readdata_from_sa) &
    ({32 {~(clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port & clock_crossing_bridge_m1_read)}} | touchPanel_spi_spi_control_port_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign clock_crossing_bridge_m1_waitrequest = ~clock_crossing_bridge_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_latency_counter <= 0;
      else 
        clock_crossing_bridge_m1_latency_counter <= p1_clock_crossing_bridge_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_clock_crossing_bridge_m1_latency_counter = ((clock_crossing_bridge_m1_run & clock_crossing_bridge_m1_read))? latency_load_value :
    (clock_crossing_bridge_m1_latency_counter)? clock_crossing_bridge_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //clock_crossing_bridge_m1_reset_n assignment, which is an e_assign
  assign clock_crossing_bridge_m1_reset_n = reset_n;

  //mux clock_crossing_bridge_m1_endofpacket, which is an e_mux
  assign clock_crossing_bridge_m1_endofpacket = touchPanel_spi_spi_control_port_endofpacket_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clock_crossing_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_address_last_time <= 0;
      else 
        clock_crossing_bridge_m1_address_last_time <= clock_crossing_bridge_m1_address;
    end


  //clock_crossing_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= clock_crossing_bridge_m1_waitrequest & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
    end


  //clock_crossing_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_bridge_m1_address != clock_crossing_bridge_m1_address_last_time))
        begin
          $write("%0d ns: clock_crossing_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_byteenable_last_time <= 0;
      else 
        clock_crossing_bridge_m1_byteenable_last_time <= clock_crossing_bridge_m1_byteenable;
    end


  //clock_crossing_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_bridge_m1_byteenable != clock_crossing_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: clock_crossing_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_read_last_time <= 0;
      else 
        clock_crossing_bridge_m1_read_last_time <= clock_crossing_bridge_m1_read;
    end


  //clock_crossing_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_bridge_m1_read != clock_crossing_bridge_m1_read_last_time))
        begin
          $write("%0d ns: clock_crossing_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_write_last_time <= 0;
      else 
        clock_crossing_bridge_m1_write_last_time <= clock_crossing_bridge_m1_write;
    end


  //clock_crossing_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_bridge_m1_write != clock_crossing_bridge_m1_write_last_time))
        begin
          $write("%0d ns: clock_crossing_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //clock_crossing_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clock_crossing_bridge_m1_writedata_last_time <= 0;
      else 
        clock_crossing_bridge_m1_writedata_last_time <= clock_crossing_bridge_m1_writedata;
    end


  //clock_crossing_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (clock_crossing_bridge_m1_writedata != clock_crossing_bridge_m1_writedata_last_time) & clock_crossing_bridge_m1_write)
        begin
          $write("%0d ns: clock_crossing_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clock_crossing_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module colour_lookup_table_s1_arbitrator (
                                           // inputs:
                                            clk,
                                            colour_lookup_table_s1_readdata,
                                            pipeline_bridge_m1_address_to_slave,
                                            pipeline_bridge_m1_burstcount,
                                            pipeline_bridge_m1_byteenable,
                                            pipeline_bridge_m1_chipselect,
                                            pipeline_bridge_m1_latency_counter,
                                            pipeline_bridge_m1_read,
                                            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                            pipeline_bridge_m1_write,
                                            pipeline_bridge_m1_writedata,
                                            reset_n,

                                           // outputs:
                                            colour_lookup_table_s1_address,
                                            colour_lookup_table_s1_byteenable,
                                            colour_lookup_table_s1_chipselect,
                                            colour_lookup_table_s1_clken,
                                            colour_lookup_table_s1_readdata_from_sa,
                                            colour_lookup_table_s1_reset,
                                            colour_lookup_table_s1_write,
                                            colour_lookup_table_s1_writedata,
                                            d1_colour_lookup_table_s1_end_xfer,
                                            pipeline_bridge_m1_granted_colour_lookup_table_s1,
                                            pipeline_bridge_m1_qualified_request_colour_lookup_table_s1,
                                            pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1,
                                            pipeline_bridge_m1_requests_colour_lookup_table_s1
                                         )
;

  output  [  7: 0] colour_lookup_table_s1_address;
  output  [  3: 0] colour_lookup_table_s1_byteenable;
  output           colour_lookup_table_s1_chipselect;
  output           colour_lookup_table_s1_clken;
  output  [ 31: 0] colour_lookup_table_s1_readdata_from_sa;
  output           colour_lookup_table_s1_reset;
  output           colour_lookup_table_s1_write;
  output  [ 31: 0] colour_lookup_table_s1_writedata;
  output           d1_colour_lookup_table_s1_end_xfer;
  output           pipeline_bridge_m1_granted_colour_lookup_table_s1;
  output           pipeline_bridge_m1_qualified_request_colour_lookup_table_s1;
  output           pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1;
  output           pipeline_bridge_m1_requests_colour_lookup_table_s1;
  input            clk;
  input   [ 31: 0] colour_lookup_table_s1_readdata;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  wire    [  7: 0] colour_lookup_table_s1_address;
  wire             colour_lookup_table_s1_allgrants;
  wire             colour_lookup_table_s1_allow_new_arb_cycle;
  wire             colour_lookup_table_s1_any_bursting_master_saved_grant;
  wire             colour_lookup_table_s1_any_continuerequest;
  wire             colour_lookup_table_s1_arb_counter_enable;
  reg              colour_lookup_table_s1_arb_share_counter;
  wire             colour_lookup_table_s1_arb_share_counter_next_value;
  wire             colour_lookup_table_s1_arb_share_set_values;
  wire             colour_lookup_table_s1_beginbursttransfer_internal;
  wire             colour_lookup_table_s1_begins_xfer;
  wire    [  3: 0] colour_lookup_table_s1_byteenable;
  wire             colour_lookup_table_s1_chipselect;
  wire             colour_lookup_table_s1_clken;
  wire             colour_lookup_table_s1_end_xfer;
  wire             colour_lookup_table_s1_firsttransfer;
  wire             colour_lookup_table_s1_grant_vector;
  wire             colour_lookup_table_s1_in_a_read_cycle;
  wire             colour_lookup_table_s1_in_a_write_cycle;
  wire             colour_lookup_table_s1_master_qreq_vector;
  wire             colour_lookup_table_s1_non_bursting_master_requests;
  wire    [ 31: 0] colour_lookup_table_s1_readdata_from_sa;
  reg              colour_lookup_table_s1_reg_firsttransfer;
  wire             colour_lookup_table_s1_reset;
  reg              colour_lookup_table_s1_slavearbiterlockenable;
  wire             colour_lookup_table_s1_slavearbiterlockenable2;
  wire             colour_lookup_table_s1_unreg_firsttransfer;
  wire             colour_lookup_table_s1_waits_for_read;
  wire             colour_lookup_table_s1_waits_for_write;
  wire             colour_lookup_table_s1_write;
  wire    [ 31: 0] colour_lookup_table_s1_writedata;
  reg              d1_colour_lookup_table_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_colour_lookup_table_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_qualified_request_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1;
  reg              pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register;
  wire             pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register_in;
  wire             pipeline_bridge_m1_requests_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_saved_grant_colour_lookup_table_s1;
  wire    [ 26: 0] shifted_address_to_colour_lookup_table_s1_from_pipeline_bridge_m1;
  wire             wait_for_colour_lookup_table_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~colour_lookup_table_s1_end_xfer;
    end


  assign colour_lookup_table_s1_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_colour_lookup_table_s1));
  //assign colour_lookup_table_s1_readdata_from_sa = colour_lookup_table_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign colour_lookup_table_s1_readdata_from_sa = colour_lookup_table_s1_readdata;

  assign pipeline_bridge_m1_requests_colour_lookup_table_s1 = ({pipeline_bridge_m1_address_to_slave[26 : 10] , 10'b0} == 27'h4401c00) & pipeline_bridge_m1_chipselect;
  //colour_lookup_table_s1_arb_share_counter set values, which is an e_mux
  assign colour_lookup_table_s1_arb_share_set_values = 1;

  //colour_lookup_table_s1_non_bursting_master_requests mux, which is an e_mux
  assign colour_lookup_table_s1_non_bursting_master_requests = pipeline_bridge_m1_requests_colour_lookup_table_s1;

  //colour_lookup_table_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign colour_lookup_table_s1_any_bursting_master_saved_grant = 0;

  //colour_lookup_table_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign colour_lookup_table_s1_arb_share_counter_next_value = colour_lookup_table_s1_firsttransfer ? (colour_lookup_table_s1_arb_share_set_values - 1) : |colour_lookup_table_s1_arb_share_counter ? (colour_lookup_table_s1_arb_share_counter - 1) : 0;

  //colour_lookup_table_s1_allgrants all slave grants, which is an e_mux
  assign colour_lookup_table_s1_allgrants = |colour_lookup_table_s1_grant_vector;

  //colour_lookup_table_s1_end_xfer assignment, which is an e_assign
  assign colour_lookup_table_s1_end_xfer = ~(colour_lookup_table_s1_waits_for_read | colour_lookup_table_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_colour_lookup_table_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_colour_lookup_table_s1 = colour_lookup_table_s1_end_xfer & (~colour_lookup_table_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //colour_lookup_table_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign colour_lookup_table_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_colour_lookup_table_s1 & colour_lookup_table_s1_allgrants) | (end_xfer_arb_share_counter_term_colour_lookup_table_s1 & ~colour_lookup_table_s1_non_bursting_master_requests);

  //colour_lookup_table_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s1_arb_share_counter <= 0;
      else if (colour_lookup_table_s1_arb_counter_enable)
          colour_lookup_table_s1_arb_share_counter <= colour_lookup_table_s1_arb_share_counter_next_value;
    end


  //colour_lookup_table_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s1_slavearbiterlockenable <= 0;
      else if ((|colour_lookup_table_s1_master_qreq_vector & end_xfer_arb_share_counter_term_colour_lookup_table_s1) | (end_xfer_arb_share_counter_term_colour_lookup_table_s1 & ~colour_lookup_table_s1_non_bursting_master_requests))
          colour_lookup_table_s1_slavearbiterlockenable <= |colour_lookup_table_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 colour_lookup_table/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = colour_lookup_table_s1_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //colour_lookup_table_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign colour_lookup_table_s1_slavearbiterlockenable2 = |colour_lookup_table_s1_arb_share_counter_next_value;

  //pipeline_bridge/m1 colour_lookup_table/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = colour_lookup_table_s1_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //colour_lookup_table_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign colour_lookup_table_s1_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_colour_lookup_table_s1 = pipeline_bridge_m1_requests_colour_lookup_table_s1 & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((1 < pipeline_bridge_m1_latency_counter) | (|pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register))));
  //pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register_in = pipeline_bridge_m1_granted_colour_lookup_table_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~colour_lookup_table_s1_waits_for_read;

  //shift register p1 pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register = {pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register, pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register_in};

  //pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register <= 0;
      else 
        pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register <= p1_pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register;
    end


  //local readdatavalid pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1 = pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1_shift_register;

  //colour_lookup_table_s1_writedata mux, which is an e_mux
  assign colour_lookup_table_s1_writedata = pipeline_bridge_m1_writedata;

  //mux colour_lookup_table_s1_clken, which is an e_mux
  assign colour_lookup_table_s1_clken = 1'b1;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_colour_lookup_table_s1 = pipeline_bridge_m1_qualified_request_colour_lookup_table_s1;

  //pipeline_bridge/m1 saved-grant colour_lookup_table/s1, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_colour_lookup_table_s1 = pipeline_bridge_m1_requests_colour_lookup_table_s1;

  //allow new arb cycle for colour_lookup_table/s1, which is an e_assign
  assign colour_lookup_table_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign colour_lookup_table_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign colour_lookup_table_s1_master_qreq_vector = 1;

  //~colour_lookup_table_s1_reset assignment, which is an e_assign
  assign colour_lookup_table_s1_reset = ~reset_n;

  assign colour_lookup_table_s1_chipselect = pipeline_bridge_m1_granted_colour_lookup_table_s1;
  //colour_lookup_table_s1_firsttransfer first transaction, which is an e_assign
  assign colour_lookup_table_s1_firsttransfer = colour_lookup_table_s1_begins_xfer ? colour_lookup_table_s1_unreg_firsttransfer : colour_lookup_table_s1_reg_firsttransfer;

  //colour_lookup_table_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign colour_lookup_table_s1_unreg_firsttransfer = ~(colour_lookup_table_s1_slavearbiterlockenable & colour_lookup_table_s1_any_continuerequest);

  //colour_lookup_table_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s1_reg_firsttransfer <= 1'b1;
      else if (colour_lookup_table_s1_begins_xfer)
          colour_lookup_table_s1_reg_firsttransfer <= colour_lookup_table_s1_unreg_firsttransfer;
    end


  //colour_lookup_table_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign colour_lookup_table_s1_beginbursttransfer_internal = colour_lookup_table_s1_begins_xfer;

  //colour_lookup_table_s1_write assignment, which is an e_mux
  assign colour_lookup_table_s1_write = pipeline_bridge_m1_granted_colour_lookup_table_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_colour_lookup_table_s1_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //colour_lookup_table_s1_address mux, which is an e_mux
  assign colour_lookup_table_s1_address = shifted_address_to_colour_lookup_table_s1_from_pipeline_bridge_m1 >> 2;

  //d1_colour_lookup_table_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_colour_lookup_table_s1_end_xfer <= 1;
      else 
        d1_colour_lookup_table_s1_end_xfer <= colour_lookup_table_s1_end_xfer;
    end


  //colour_lookup_table_s1_waits_for_read in a cycle, which is an e_mux
  assign colour_lookup_table_s1_waits_for_read = colour_lookup_table_s1_in_a_read_cycle & 0;

  //colour_lookup_table_s1_in_a_read_cycle assignment, which is an e_assign
  assign colour_lookup_table_s1_in_a_read_cycle = pipeline_bridge_m1_granted_colour_lookup_table_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = colour_lookup_table_s1_in_a_read_cycle;

  //colour_lookup_table_s1_waits_for_write in a cycle, which is an e_mux
  assign colour_lookup_table_s1_waits_for_write = colour_lookup_table_s1_in_a_write_cycle & 0;

  //colour_lookup_table_s1_in_a_write_cycle assignment, which is an e_assign
  assign colour_lookup_table_s1_in_a_write_cycle = pipeline_bridge_m1_granted_colour_lookup_table_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = colour_lookup_table_s1_in_a_write_cycle;

  assign wait_for_colour_lookup_table_s1_counter = 0;
  //colour_lookup_table_s1_byteenable byte enable port mux, which is an e_mux
  assign colour_lookup_table_s1_byteenable = (pipeline_bridge_m1_granted_colour_lookup_table_s1)? pipeline_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //colour_lookup_table/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_colour_lookup_table_s1 && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave colour_lookup_table/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module colour_lookup_table_s2_arbitrator (
                                           // inputs:
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave,
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported,
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter,
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read,
                                            clk,
                                            colour_lookup_table_s2_readdata,
                                            dummy_master_inst_m0_address_to_slave,
                                            dummy_master_inst_m0_write,
                                            dummy_master_inst_m0_writedata,
                                            reset_n,

                                           // outputs:
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2,
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2,
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2,
                                            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2,
                                            colour_lookup_table_s2_address,
                                            colour_lookup_table_s2_byteenable,
                                            colour_lookup_table_s2_chipselect,
                                            colour_lookup_table_s2_clken,
                                            colour_lookup_table_s2_readdata_from_sa,
                                            colour_lookup_table_s2_reset,
                                            colour_lookup_table_s2_write,
                                            colour_lookup_table_s2_writedata,
                                            d1_colour_lookup_table_s2_end_xfer,
                                            dummy_master_inst_granted_colour_lookup_table_s2,
                                            dummy_master_inst_qualified_request_colour_lookup_table_s2,
                                            dummy_master_inst_requests_colour_lookup_table_s2
                                         )
;

  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2;
  output  [  7: 0] colour_lookup_table_s2_address;
  output  [  3: 0] colour_lookup_table_s2_byteenable;
  output           colour_lookup_table_s2_chipselect;
  output           colour_lookup_table_s2_clken;
  output  [ 31: 0] colour_lookup_table_s2_readdata_from_sa;
  output           colour_lookup_table_s2_reset;
  output           colour_lookup_table_s2_write;
  output  [ 31: 0] colour_lookup_table_s2_writedata;
  output           d1_colour_lookup_table_s2_end_xfer;
  output           dummy_master_inst_granted_colour_lookup_table_s2;
  output           dummy_master_inst_qualified_request_colour_lookup_table_s2;
  output           dummy_master_inst_requests_colour_lookup_table_s2;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read;
  input            clk;
  input   [ 31: 0] colour_lookup_table_s2_readdata;
  input   [ 31: 0] dummy_master_inst_m0_address_to_slave;
  input            dummy_master_inst_m0_write;
  input   [ 31: 0] dummy_master_inst_m0_writedata;
  input            reset_n;

  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbiterlock;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbiterlock2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2;
  reg              accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register_in;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_saved_grant_colour_lookup_table_s2;
  wire    [  7: 0] colour_lookup_table_s2_address;
  wire             colour_lookup_table_s2_allgrants;
  wire             colour_lookup_table_s2_allow_new_arb_cycle;
  wire             colour_lookup_table_s2_any_bursting_master_saved_grant;
  wire             colour_lookup_table_s2_any_continuerequest;
  reg     [  1: 0] colour_lookup_table_s2_arb_addend;
  wire             colour_lookup_table_s2_arb_counter_enable;
  reg              colour_lookup_table_s2_arb_share_counter;
  wire             colour_lookup_table_s2_arb_share_counter_next_value;
  wire             colour_lookup_table_s2_arb_share_set_values;
  wire    [  1: 0] colour_lookup_table_s2_arb_winner;
  wire             colour_lookup_table_s2_arbitration_holdoff_internal;
  wire             colour_lookup_table_s2_beginbursttransfer_internal;
  wire             colour_lookup_table_s2_begins_xfer;
  wire    [  3: 0] colour_lookup_table_s2_byteenable;
  wire             colour_lookup_table_s2_chipselect;
  wire    [  3: 0] colour_lookup_table_s2_chosen_master_double_vector;
  wire    [  1: 0] colour_lookup_table_s2_chosen_master_rot_left;
  wire             colour_lookup_table_s2_clken;
  wire             colour_lookup_table_s2_end_xfer;
  wire             colour_lookup_table_s2_firsttransfer;
  wire    [  1: 0] colour_lookup_table_s2_grant_vector;
  wire             colour_lookup_table_s2_in_a_read_cycle;
  wire             colour_lookup_table_s2_in_a_write_cycle;
  wire    [  1: 0] colour_lookup_table_s2_master_qreq_vector;
  wire             colour_lookup_table_s2_non_bursting_master_requests;
  wire    [ 31: 0] colour_lookup_table_s2_readdata_from_sa;
  reg              colour_lookup_table_s2_reg_firsttransfer;
  wire             colour_lookup_table_s2_reset;
  reg     [  1: 0] colour_lookup_table_s2_saved_chosen_master_vector;
  reg              colour_lookup_table_s2_slavearbiterlockenable;
  wire             colour_lookup_table_s2_slavearbiterlockenable2;
  wire             colour_lookup_table_s2_unreg_firsttransfer;
  wire             colour_lookup_table_s2_waits_for_read;
  wire             colour_lookup_table_s2_waits_for_write;
  wire             colour_lookup_table_s2_write;
  wire    [ 31: 0] colour_lookup_table_s2_writedata;
  reg              d1_colour_lookup_table_s2_end_xfer;
  reg              d1_reasons_to_wait;
  wire             dummy_master_inst_granted_colour_lookup_table_s2;
  wire             dummy_master_inst_m0_arbiterlock;
  wire             dummy_master_inst_m0_arbiterlock2;
  wire             dummy_master_inst_m0_continuerequest;
  wire             dummy_master_inst_qualified_request_colour_lookup_table_s2;
  wire             dummy_master_inst_requests_colour_lookup_table_s2;
  wire             dummy_master_inst_saved_grant_colour_lookup_table_s2;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_colour_lookup_table_s2;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_slave_colour_lookup_table_s2;
  reg              last_cycle_dummy_master_inst_m0_granted_slave_colour_lookup_table_s2;
  wire             p1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register;
  wire    [ 31: 0] shifted_address_to_colour_lookup_table_s2_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0;
  wire    [ 31: 0] shifted_address_to_colour_lookup_table_s2_from_dummy_master_inst_m0;
  wire             wait_for_colour_lookup_table_s2_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~colour_lookup_table_s2_end_xfer;
    end


  assign colour_lookup_table_s2_begins_xfer = ~d1_reasons_to_wait & ((accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2 | dummy_master_inst_qualified_request_colour_lookup_table_s2));
  //assign colour_lookup_table_s2_readdata_from_sa = colour_lookup_table_s2_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign colour_lookup_table_s2_readdata_from_sa = colour_lookup_table_s2_readdata;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2 = (({accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave[31 : 10] , 10'b0} == 32'h4401c00) & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read)) & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read;
  //colour_lookup_table_s2_arb_share_counter set values, which is an e_mux
  assign colour_lookup_table_s2_arb_share_set_values = 1;

  //colour_lookup_table_s2_non_bursting_master_requests mux, which is an e_mux
  assign colour_lookup_table_s2_non_bursting_master_requests = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2 |
    dummy_master_inst_requests_colour_lookup_table_s2 |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2 |
    dummy_master_inst_requests_colour_lookup_table_s2;

  //colour_lookup_table_s2_any_bursting_master_saved_grant mux, which is an e_mux
  assign colour_lookup_table_s2_any_bursting_master_saved_grant = 0;

  //colour_lookup_table_s2_arb_share_counter_next_value assignment, which is an e_assign
  assign colour_lookup_table_s2_arb_share_counter_next_value = colour_lookup_table_s2_firsttransfer ? (colour_lookup_table_s2_arb_share_set_values - 1) : |colour_lookup_table_s2_arb_share_counter ? (colour_lookup_table_s2_arb_share_counter - 1) : 0;

  //colour_lookup_table_s2_allgrants all slave grants, which is an e_mux
  assign colour_lookup_table_s2_allgrants = (|colour_lookup_table_s2_grant_vector) |
    (|colour_lookup_table_s2_grant_vector) |
    (|colour_lookup_table_s2_grant_vector) |
    (|colour_lookup_table_s2_grant_vector);

  //colour_lookup_table_s2_end_xfer assignment, which is an e_assign
  assign colour_lookup_table_s2_end_xfer = ~(colour_lookup_table_s2_waits_for_read | colour_lookup_table_s2_waits_for_write);

  //end_xfer_arb_share_counter_term_colour_lookup_table_s2 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_colour_lookup_table_s2 = colour_lookup_table_s2_end_xfer & (~colour_lookup_table_s2_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //colour_lookup_table_s2_arb_share_counter arbitration counter enable, which is an e_assign
  assign colour_lookup_table_s2_arb_counter_enable = (end_xfer_arb_share_counter_term_colour_lookup_table_s2 & colour_lookup_table_s2_allgrants) | (end_xfer_arb_share_counter_term_colour_lookup_table_s2 & ~colour_lookup_table_s2_non_bursting_master_requests);

  //colour_lookup_table_s2_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s2_arb_share_counter <= 0;
      else if (colour_lookup_table_s2_arb_counter_enable)
          colour_lookup_table_s2_arb_share_counter <= colour_lookup_table_s2_arb_share_counter_next_value;
    end


  //colour_lookup_table_s2_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s2_slavearbiterlockenable <= 0;
      else if ((|colour_lookup_table_s2_master_qreq_vector & end_xfer_arb_share_counter_term_colour_lookup_table_s2) | (end_xfer_arb_share_counter_term_colour_lookup_table_s2 & ~colour_lookup_table_s2_non_bursting_master_requests))
          colour_lookup_table_s2_slavearbiterlockenable <= |colour_lookup_table_s2_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 colour_lookup_table/s2 arbiterlock, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbiterlock = colour_lookup_table_s2_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_continuerequest;

  //colour_lookup_table_s2_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign colour_lookup_table_s2_slavearbiterlockenable2 = |colour_lookup_table_s2_arb_share_counter_next_value;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 colour_lookup_table/s2 arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbiterlock2 = colour_lookup_table_s2_slavearbiterlockenable2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_continuerequest;

  //dummy_master_inst/m0 colour_lookup_table/s2 arbiterlock, which is an e_assign
  assign dummy_master_inst_m0_arbiterlock = colour_lookup_table_s2_slavearbiterlockenable & dummy_master_inst_m0_continuerequest;

  //dummy_master_inst/m0 colour_lookup_table/s2 arbiterlock2, which is an e_assign
  assign dummy_master_inst_m0_arbiterlock2 = colour_lookup_table_s2_slavearbiterlockenable2 & dummy_master_inst_m0_continuerequest;

  //dummy_master_inst/m0 granted colour_lookup_table/s2 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_dummy_master_inst_m0_granted_slave_colour_lookup_table_s2 <= 0;
      else 
        last_cycle_dummy_master_inst_m0_granted_slave_colour_lookup_table_s2 <= dummy_master_inst_saved_grant_colour_lookup_table_s2 ? 1 : (colour_lookup_table_s2_arbitration_holdoff_internal | ~dummy_master_inst_requests_colour_lookup_table_s2) ? 0 : last_cycle_dummy_master_inst_m0_granted_slave_colour_lookup_table_s2;
    end


  //dummy_master_inst_m0_continuerequest continued request, which is an e_mux
  assign dummy_master_inst_m0_continuerequest = last_cycle_dummy_master_inst_m0_granted_slave_colour_lookup_table_s2 & dummy_master_inst_requests_colour_lookup_table_s2;

  //colour_lookup_table_s2_any_continuerequest at least one master continues requesting, which is an e_mux
  assign colour_lookup_table_s2_any_continuerequest = dummy_master_inst_m0_continuerequest |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_continuerequest;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2 & ~(dummy_master_inst_m0_arbiterlock);
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register_in mux for readlatency shift register, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register_in = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read & ~colour_lookup_table_s2_waits_for_read;

  //shift register p1 accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported)? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register_in :
    {accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register, accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register_in};

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register <= 0;
      else 
        accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register <= p1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register;
    end


  //local readdatavalid accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2_shift_register;

  //mux colour_lookup_table_s2_clken, which is an e_mux
  assign colour_lookup_table_s2_clken = 1'b1;

  assign dummy_master_inst_requests_colour_lookup_table_s2 = (({dummy_master_inst_m0_address_to_slave[31 : 10] , 10'b0} == 32'h4401c00) & (dummy_master_inst_m0_write)) & dummy_master_inst_m0_write;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 granted colour_lookup_table/s2 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_slave_colour_lookup_table_s2 <= 0;
      else 
        last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_slave_colour_lookup_table_s2 <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_saved_grant_colour_lookup_table_s2 ? 1 : (colour_lookup_table_s2_arbitration_holdoff_internal | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2) ? 0 : last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_slave_colour_lookup_table_s2;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_continuerequest continued request, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_continuerequest = last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_slave_colour_lookup_table_s2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2;

  assign dummy_master_inst_qualified_request_colour_lookup_table_s2 = dummy_master_inst_requests_colour_lookup_table_s2 & ~(accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbiterlock);
  //colour_lookup_table_s2_writedata mux, which is an e_mux
  assign colour_lookup_table_s2_writedata = dummy_master_inst_m0_writedata;

  //allow new arb cycle for colour_lookup_table/s2, which is an e_assign
  assign colour_lookup_table_s2_allow_new_arb_cycle = ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbiterlock & ~dummy_master_inst_m0_arbiterlock;

  //dummy_master_inst/m0 assignment into master qualified-requests vector for colour_lookup_table/s2, which is an e_assign
  assign colour_lookup_table_s2_master_qreq_vector[0] = dummy_master_inst_qualified_request_colour_lookup_table_s2;

  //dummy_master_inst/m0 grant colour_lookup_table/s2, which is an e_assign
  assign dummy_master_inst_granted_colour_lookup_table_s2 = colour_lookup_table_s2_grant_vector[0];

  //dummy_master_inst/m0 saved-grant colour_lookup_table/s2, which is an e_assign
  assign dummy_master_inst_saved_grant_colour_lookup_table_s2 = colour_lookup_table_s2_arb_winner[0] && dummy_master_inst_requests_colour_lookup_table_s2;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 assignment into master qualified-requests vector for colour_lookup_table/s2, which is an e_assign
  assign colour_lookup_table_s2_master_qreq_vector[1] = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 grant colour_lookup_table/s2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2 = colour_lookup_table_s2_grant_vector[1];

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 saved-grant colour_lookup_table/s2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_saved_grant_colour_lookup_table_s2 = colour_lookup_table_s2_arb_winner[1] && accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2;

  //colour_lookup_table/s2 chosen-master double-vector, which is an e_assign
  assign colour_lookup_table_s2_chosen_master_double_vector = {colour_lookup_table_s2_master_qreq_vector, colour_lookup_table_s2_master_qreq_vector} & ({~colour_lookup_table_s2_master_qreq_vector, ~colour_lookup_table_s2_master_qreq_vector} + colour_lookup_table_s2_arb_addend);

  //stable onehot encoding of arb winner
  assign colour_lookup_table_s2_arb_winner = (colour_lookup_table_s2_allow_new_arb_cycle & | colour_lookup_table_s2_grant_vector) ? colour_lookup_table_s2_grant_vector : colour_lookup_table_s2_saved_chosen_master_vector;

  //saved colour_lookup_table_s2_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s2_saved_chosen_master_vector <= 0;
      else if (colour_lookup_table_s2_allow_new_arb_cycle)
          colour_lookup_table_s2_saved_chosen_master_vector <= |colour_lookup_table_s2_grant_vector ? colour_lookup_table_s2_grant_vector : colour_lookup_table_s2_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign colour_lookup_table_s2_grant_vector = {(colour_lookup_table_s2_chosen_master_double_vector[1] | colour_lookup_table_s2_chosen_master_double_vector[3]),
    (colour_lookup_table_s2_chosen_master_double_vector[0] | colour_lookup_table_s2_chosen_master_double_vector[2])};

  //colour_lookup_table/s2 chosen master rotated left, which is an e_assign
  assign colour_lookup_table_s2_chosen_master_rot_left = (colour_lookup_table_s2_arb_winner << 1) ? (colour_lookup_table_s2_arb_winner << 1) : 1;

  //colour_lookup_table/s2's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s2_arb_addend <= 1;
      else if (|colour_lookup_table_s2_grant_vector)
          colour_lookup_table_s2_arb_addend <= colour_lookup_table_s2_end_xfer? colour_lookup_table_s2_chosen_master_rot_left : colour_lookup_table_s2_grant_vector;
    end


  //~colour_lookup_table_s2_reset assignment, which is an e_assign
  assign colour_lookup_table_s2_reset = ~reset_n;

  assign colour_lookup_table_s2_chipselect = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2 | dummy_master_inst_granted_colour_lookup_table_s2;
  //colour_lookup_table_s2_firsttransfer first transaction, which is an e_assign
  assign colour_lookup_table_s2_firsttransfer = colour_lookup_table_s2_begins_xfer ? colour_lookup_table_s2_unreg_firsttransfer : colour_lookup_table_s2_reg_firsttransfer;

  //colour_lookup_table_s2_unreg_firsttransfer first transaction, which is an e_assign
  assign colour_lookup_table_s2_unreg_firsttransfer = ~(colour_lookup_table_s2_slavearbiterlockenable & colour_lookup_table_s2_any_continuerequest);

  //colour_lookup_table_s2_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          colour_lookup_table_s2_reg_firsttransfer <= 1'b1;
      else if (colour_lookup_table_s2_begins_xfer)
          colour_lookup_table_s2_reg_firsttransfer <= colour_lookup_table_s2_unreg_firsttransfer;
    end


  //colour_lookup_table_s2_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign colour_lookup_table_s2_beginbursttransfer_internal = colour_lookup_table_s2_begins_xfer;

  //colour_lookup_table_s2_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign colour_lookup_table_s2_arbitration_holdoff_internal = colour_lookup_table_s2_begins_xfer & colour_lookup_table_s2_firsttransfer;

  //colour_lookup_table_s2_write assignment, which is an e_mux
  assign colour_lookup_table_s2_write = dummy_master_inst_granted_colour_lookup_table_s2 & dummy_master_inst_m0_write;

  assign shifted_address_to_colour_lookup_table_s2_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave;
  //colour_lookup_table_s2_address mux, which is an e_mux
  assign colour_lookup_table_s2_address = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2)? (shifted_address_to_colour_lookup_table_s2_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0 >> 2) :
    (shifted_address_to_colour_lookup_table_s2_from_dummy_master_inst_m0 >> 2);

  assign shifted_address_to_colour_lookup_table_s2_from_dummy_master_inst_m0 = dummy_master_inst_m0_address_to_slave;
  //d1_colour_lookup_table_s2_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_colour_lookup_table_s2_end_xfer <= 1;
      else 
        d1_colour_lookup_table_s2_end_xfer <= colour_lookup_table_s2_end_xfer;
    end


  //colour_lookup_table_s2_waits_for_read in a cycle, which is an e_mux
  assign colour_lookup_table_s2_waits_for_read = colour_lookup_table_s2_in_a_read_cycle & 0;

  //colour_lookup_table_s2_in_a_read_cycle assignment, which is an e_assign
  assign colour_lookup_table_s2_in_a_read_cycle = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = colour_lookup_table_s2_in_a_read_cycle;

  //colour_lookup_table_s2_waits_for_write in a cycle, which is an e_mux
  assign colour_lookup_table_s2_waits_for_write = colour_lookup_table_s2_in_a_write_cycle & 0;

  //colour_lookup_table_s2_in_a_write_cycle assignment, which is an e_assign
  assign colour_lookup_table_s2_in_a_write_cycle = dummy_master_inst_granted_colour_lookup_table_s2 & dummy_master_inst_m0_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = colour_lookup_table_s2_in_a_write_cycle;

  assign wait_for_colour_lookup_table_s2_counter = 0;
  //colour_lookup_table_s2_byteenable byte enable port mux, which is an e_mux
  assign colour_lookup_table_s2_byteenable = (dummy_master_inst_granted_colour_lookup_table_s2)? {4 {1'b1}} :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //colour_lookup_table/s2 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2 + dummy_master_inst_granted_colour_lookup_table_s2 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_saved_grant_colour_lookup_table_s2 + dummy_master_inst_saved_grant_colour_lookup_table_s2 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           pipeline_bridge_m1_address_to_slave,
                                           pipeline_bridge_m1_burstcount,
                                           pipeline_bridge_m1_byteenable,
                                           pipeline_bridge_m1_chipselect,
                                           pipeline_bridge_m1_debugaccess,
                                           pipeline_bridge_m1_latency_counter,
                                           pipeline_bridge_m1_read,
                                           pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                           pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                           pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                           pipeline_bridge_m1_write,
                                           pipeline_bridge_m1_writedata,
                                           reset_n,

                                          // outputs:
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer,
                                           pipeline_bridge_m1_granted_cpu_jtag_debug_module,
                                           pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module,
                                           pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module,
                                           pipeline_bridge_m1_requests_cpu_jtag_debug_module
                                        )
;

  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  output           pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  output           pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  output           pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  output           pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  input            clk;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_debugaccess;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg              cpu_jtag_debug_module_arb_share_counter;
  wire             cpu_jtag_debug_module_arb_share_counter_next_value;
  wire             cpu_jtag_debug_module_arb_share_set_values;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire             cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire             cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_saved_grant_cpu_jtag_debug_module;
  wire    [ 26: 0] shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign pipeline_bridge_m1_requests_cpu_jtag_debug_module = ({pipeline_bridge_m1_address_to_slave[26 : 11] , 11'b0} == 27'h4401000) & pipeline_bridge_m1_chipselect;
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = 1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = pipeline_bridge_m1_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = |cpu_jtag_debug_module_grant_vector;

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //pipeline_bridge/m1 cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_assign
  assign cpu_jtag_debug_module_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module = pipeline_bridge_m1_requests_cpu_jtag_debug_module & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0) | (|pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~cpu_jtag_debug_module_waits_for_read;

  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = pipeline_bridge_m1_writedata;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_cpu_jtag_debug_module = pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;

  //pipeline_bridge/m1 saved-grant cpu/jtag_debug_module, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_cpu_jtag_debug_module = pipeline_bridge_m1_requests_cpu_jtag_debug_module;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign cpu_jtag_debug_module_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign cpu_jtag_debug_module_master_qreq_vector = 1;

  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1 >> 2;

  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (pipeline_bridge_m1_granted_cpu_jtag_debug_module)? pipeline_bridge_m1_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (pipeline_bridge_m1_granted_cpu_jtag_debug_module)? pipeline_bridge_m1_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_cpu_jtag_debug_module && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                                       // inputs:
                                                                                        clk,
                                                                                        data_in,
                                                                                        reset_n,

                                                                                       // outputs:
                                                                                        data_out
                                                                                     )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module push_buttons_s1_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                           // inputs:
                                                                            clk,
                                                                            data_in,
                                                                            reset_n,

                                                                           // outputs:
                                                                            data_out
                                                                         )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_tick_s1_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                          // inputs:
                                                                           clk,
                                                                           data_in,
                                                                           reset_n,

                                                                          // outputs:
                                                                           data_out
                                                                        )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module touchPanel_irq_n_s1_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                               // inputs:
                                                                                clk,
                                                                                data_in,
                                                                                reset_n,

                                                                               // outputs:
                                                                                data_out
                                                                             )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module touchPanel_spi_spi_control_port_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                                           // inputs:
                                                                                            clk,
                                                                                            data_in,
                                                                                            reset_n,

                                                                                           // outputs:
                                                                                            data_out
                                                                                         )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa,
                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa,
                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa,
                                     clk,
                                     cpu_data_master_address,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                     cpu_data_master_granted_pipeline_bridge_s1,
                                     cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                     cpu_data_master_qualified_request_pipeline_bridge_s1,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                     cpu_data_master_read_data_valid_pipeline_bridge_s1,
                                     cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
                                     cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0,
                                     cpu_data_master_requests_pipeline_bridge_s1,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer,
                                     d1_pipeline_bridge_s1_end_xfer,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     lcd_sgdma_csr_irq_from_sa,
                                     pipeline_bridge_s1_readdata_from_sa,
                                     pipeline_bridge_s1_waitrequest_from_sa,
                                     push_buttons_s1_irq_from_sa,
                                     reset_n,
                                     system_clk,
                                     system_clk_reset_n,
                                     system_tick_s1_irq_from_sa,
                                     touchPanel_irq_n_s1_irq_from_sa,
                                     touchPanel_spi_spi_control_port_irq_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_irq,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_readdata,
                                     cpu_data_master_readdatavalid,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 27: 0] cpu_data_master_address_to_slave;
  output  [ 31: 0] cpu_data_master_irq;
  output           cpu_data_master_latency_counter;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_readdatavalid;
  output           cpu_data_master_waitrequest;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa;
  input            clk;
  input   [ 27: 0] cpu_data_master_address;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  input            cpu_data_master_granted_pipeline_bridge_s1;
  input            cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  input            cpu_data_master_qualified_request_pipeline_bridge_s1;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  input            cpu_data_master_read_data_valid_pipeline_bridge_s1;
  input            cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register;
  input            cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  input            cpu_data_master_requests_pipeline_bridge_s1;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
  input            d1_pipeline_bridge_s1_end_xfer;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input            lcd_sgdma_csr_irq_from_sa;
  input   [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  input            pipeline_bridge_s1_waitrequest_from_sa;
  input            push_buttons_s1_irq_from_sa;
  input            reset_n;
  input            system_clk;
  input            system_clk_reset_n;
  input            system_tick_s1_irq_from_sa;
  input            touchPanel_irq_n_s1_irq_from_sa;
  input            touchPanel_spi_spi_control_port_irq_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 27: 0] cpu_data_master_address_last_time;
  wire    [ 27: 0] cpu_data_master_address_to_slave;
  reg     [  3: 0] cpu_data_master_byteenable_last_time;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_is_granted_some_slave;
  reg              cpu_data_master_latency_counter;
  reg              cpu_data_master_read_but_no_slave_selected;
  reg              cpu_data_master_read_last_time;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_run;
  wire             cpu_data_master_waitrequest;
  reg              cpu_data_master_write_last_time;
  reg     [ 31: 0] cpu_data_master_writedata_last_time;
  wire             latency_load_value;
  wire             p1_cpu_data_master_latency_counter;
  wire             pre_flush_cpu_data_master_readdatavalid;
  wire             r_0;
  wire             r_2;
  wire             system_clk_jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             system_clk_push_buttons_s1_irq_from_sa;
  wire             system_clk_system_tick_s1_irq_from_sa;
  wire             system_clk_touchPanel_irq_n_s1_irq_from_sa;
  wire             system_clk_touchPanel_spi_spi_control_port_irq_from_sa;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 | ~cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0) & ((~cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0 & r_2;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_data_master_qualified_request_pipeline_bridge_s1 | ~cpu_data_master_requests_pipeline_bridge_s1) & (cpu_data_master_granted_pipeline_bridge_s1 | ~cpu_data_master_qualified_request_pipeline_bridge_s1) & ((~cpu_data_master_qualified_request_pipeline_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_pipeline_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = cpu_data_master_address[27 : 0];

  //cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_data_master_read_but_no_slave_selected <= cpu_data_master_read & cpu_data_master_run & ~cpu_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_data_master_is_granted_some_slave = cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 |
    cpu_data_master_granted_pipeline_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_data_master_readdatavalid = cpu_data_master_read_data_valid_pipeline_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_data_master_readdatavalid = cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid;

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~(cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 & cpu_data_master_read)}} | accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_pipeline_bridge_s1}} | pipeline_bridge_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_data_master_waitrequest = ~cpu_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_latency_counter <= 0;
      else 
        cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_data_master_latency_counter = ((cpu_data_master_run & cpu_data_master_read))? latency_load_value :
    (cpu_data_master_latency_counter)? cpu_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa,
    system_clk_touchPanel_irq_n_s1_irq_from_sa,
    system_clk_touchPanel_spi_spi_control_port_irq_from_sa,
    lcd_sgdma_csr_irq_from_sa,
    system_clk_system_tick_s1_irq_from_sa,
    system_clk_push_buttons_s1_irq_from_sa,
    system_clk_jtag_uart_avalon_jtag_slave_irq_from_sa};

  //jtag_uart_avalon_jtag_slave_irq_from_sa from slow_clk to system_clk
  jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_data_master_module jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (system_clk),
      .data_in  (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .data_out (system_clk_jtag_uart_avalon_jtag_slave_irq_from_sa),
      .reset_n  (system_clk_reset_n)
    );

  //push_buttons_s1_irq_from_sa from slow_clk to system_clk
  push_buttons_s1_irq_from_sa_clock_crossing_cpu_data_master_module push_buttons_s1_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (system_clk),
      .data_in  (push_buttons_s1_irq_from_sa),
      .data_out (system_clk_push_buttons_s1_irq_from_sa),
      .reset_n  (system_clk_reset_n)
    );

  //system_tick_s1_irq_from_sa from slow_clk to system_clk
  system_tick_s1_irq_from_sa_clock_crossing_cpu_data_master_module system_tick_s1_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (system_clk),
      .data_in  (system_tick_s1_irq_from_sa),
      .data_out (system_clk_system_tick_s1_irq_from_sa),
      .reset_n  (system_clk_reset_n)
    );

  //touchPanel_irq_n_s1_irq_from_sa from slow_clk to system_clk
  touchPanel_irq_n_s1_irq_from_sa_clock_crossing_cpu_data_master_module touchPanel_irq_n_s1_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (system_clk),
      .data_in  (touchPanel_irq_n_s1_irq_from_sa),
      .data_out (system_clk_touchPanel_irq_n_s1_irq_from_sa),
      .reset_n  (system_clk_reset_n)
    );

  //touchPanel_spi_spi_control_port_irq_from_sa from slow_clk to system_clk
  touchPanel_spi_spi_control_port_irq_from_sa_clock_crossing_cpu_data_master_module touchPanel_spi_spi_control_port_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (system_clk),
      .data_in  (touchPanel_spi_spi_control_port_irq_from_sa),
      .data_out (system_clk_touchPanel_spi_spi_control_port_irq_from_sa),
      .reset_n  (system_clk_reset_n)
    );


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_address_last_time <= 0;
      else 
        cpu_data_master_address_last_time <= cpu_data_master_address;
    end


  //cpu/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_data_master_waitrequest & (cpu_data_master_read | cpu_data_master_write);
    end


  //cpu_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_address != cpu_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_byteenable_last_time <= 0;
      else 
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
    end


  //cpu_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_byteenable != cpu_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_last_time <= 0;
      else 
        cpu_data_master_read_last_time <= cpu_data_master_read;
    end


  //cpu_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_read != cpu_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_write_last_time <= 0;
      else 
        cpu_data_master_write_last_time <= cpu_data_master_write;
    end


  //cpu_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_write != cpu_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_writedata_last_time <= 0;
      else 
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
    end


  //cpu_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_writedata != cpu_data_master_writedata_last_time) & cpu_data_master_write)
        begin
          $write("%0d ns: cpu_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_granted_pipeline_bridge_s1,
                                            cpu_instruction_master_qualified_request_pipeline_bridge_s1,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_pipeline_bridge_s1,
                                            cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register,
                                            cpu_instruction_master_requests_pipeline_bridge_s1,
                                            d1_pipeline_bridge_s1_end_xfer,
                                            pipeline_bridge_s1_readdata_from_sa,
                                            pipeline_bridge_s1_waitrequest_from_sa,
                                            reset_n,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 26: 0] cpu_instruction_master_address_to_slave;
  output           cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 26: 0] cpu_instruction_master_address;
  input            cpu_instruction_master_granted_pipeline_bridge_s1;
  input            cpu_instruction_master_qualified_request_pipeline_bridge_s1;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_pipeline_bridge_s1;
  input            cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register;
  input            cpu_instruction_master_requests_pipeline_bridge_s1;
  input            d1_pipeline_bridge_s1_end_xfer;
  input   [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  input            pipeline_bridge_s1_waitrequest_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] cpu_instruction_master_address_last_time;
  wire    [ 26: 0] cpu_instruction_master_address_to_slave;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg              cpu_instruction_master_latency_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             latency_load_value;
  wire             p1_cpu_instruction_master_latency_counter;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_2;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_instruction_master_qualified_request_pipeline_bridge_s1 | ~cpu_instruction_master_requests_pipeline_bridge_s1) & (cpu_instruction_master_granted_pipeline_bridge_s1 | ~cpu_instruction_master_qualified_request_pipeline_bridge_s1) & ((~cpu_instruction_master_qualified_request_pipeline_bridge_s1 | ~(cpu_instruction_master_read) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (cpu_instruction_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = cpu_instruction_master_address[26 : 0];

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_pipeline_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_pipeline_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = pipeline_bridge_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else 
        cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else 
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else 
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_frame_buffer_pipeline_bridge_m1_to_ddr_sdram_clock_crossing_bridge_s1_module (
                                                                                                   // inputs:
                                                                                                    clear_fifo,
                                                                                                    clk,
                                                                                                    data_in,
                                                                                                    read,
                                                                                                    reset_n,
                                                                                                    sync_reset,
                                                                                                    write,

                                                                                                   // outputs:
                                                                                                    data_out,
                                                                                                    empty,
                                                                                                    fifo_contains_ones_n,
                                                                                                    full
                                                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  wire             full_48;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_47;
  assign empty = !full_0;
  assign full_48 = 0;
  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    0;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_clock_crossing_bridge_s1_arbitrator (
                                                       // inputs:
                                                        clk,
                                                        ddr_sdram_clock_crossing_bridge_s1_endofpacket,
                                                        ddr_sdram_clock_crossing_bridge_s1_readdata,
                                                        ddr_sdram_clock_crossing_bridge_s1_readdatavalid,
                                                        ddr_sdram_clock_crossing_bridge_s1_waitrequest,
                                                        frame_buffer_pipeline_bridge_m1_address_to_slave,
                                                        frame_buffer_pipeline_bridge_m1_burstcount,
                                                        frame_buffer_pipeline_bridge_m1_byteenable,
                                                        frame_buffer_pipeline_bridge_m1_chipselect,
                                                        frame_buffer_pipeline_bridge_m1_latency_counter,
                                                        frame_buffer_pipeline_bridge_m1_read,
                                                        frame_buffer_pipeline_bridge_m1_write,
                                                        frame_buffer_pipeline_bridge_m1_writedata,
                                                        reset_n,

                                                       // outputs:
                                                        d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer,
                                                        ddr_sdram_clock_crossing_bridge_s1_address,
                                                        ddr_sdram_clock_crossing_bridge_s1_byteenable,
                                                        ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa,
                                                        ddr_sdram_clock_crossing_bridge_s1_nativeaddress,
                                                        ddr_sdram_clock_crossing_bridge_s1_read,
                                                        ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa,
                                                        ddr_sdram_clock_crossing_bridge_s1_reset_n,
                                                        ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa,
                                                        ddr_sdram_clock_crossing_bridge_s1_write,
                                                        ddr_sdram_clock_crossing_bridge_s1_writedata,
                                                        frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1,
                                                        frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1,
                                                        frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1,
                                                        frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register,
                                                        frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1
                                                     )
;

  output           d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer;
  output  [ 22: 0] ddr_sdram_clock_crossing_bridge_s1_address;
  output  [  3: 0] ddr_sdram_clock_crossing_bridge_s1_byteenable;
  output           ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa;
  output  [ 22: 0] ddr_sdram_clock_crossing_bridge_s1_nativeaddress;
  output           ddr_sdram_clock_crossing_bridge_s1_read;
  output  [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa;
  output           ddr_sdram_clock_crossing_bridge_s1_reset_n;
  output           ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa;
  output           ddr_sdram_clock_crossing_bridge_s1_write;
  output  [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_writedata;
  output           frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1;
  output           frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1;
  output           frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1;
  output           frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register;
  output           frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1;
  input            clk;
  input            ddr_sdram_clock_crossing_bridge_s1_endofpacket;
  input   [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_readdata;
  input            ddr_sdram_clock_crossing_bridge_s1_readdatavalid;
  input            ddr_sdram_clock_crossing_bridge_s1_waitrequest;
  input   [ 24: 0] frame_buffer_pipeline_bridge_m1_address_to_slave;
  input            frame_buffer_pipeline_bridge_m1_burstcount;
  input   [  3: 0] frame_buffer_pipeline_bridge_m1_byteenable;
  input            frame_buffer_pipeline_bridge_m1_chipselect;
  input            frame_buffer_pipeline_bridge_m1_latency_counter;
  input            frame_buffer_pipeline_bridge_m1_read;
  input            frame_buffer_pipeline_bridge_m1_write;
  input   [ 31: 0] frame_buffer_pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [ 22: 0] ddr_sdram_clock_crossing_bridge_s1_address;
  wire             ddr_sdram_clock_crossing_bridge_s1_allgrants;
  wire             ddr_sdram_clock_crossing_bridge_s1_allow_new_arb_cycle;
  wire             ddr_sdram_clock_crossing_bridge_s1_any_bursting_master_saved_grant;
  wire             ddr_sdram_clock_crossing_bridge_s1_any_continuerequest;
  wire             ddr_sdram_clock_crossing_bridge_s1_arb_counter_enable;
  reg              ddr_sdram_clock_crossing_bridge_s1_arb_share_counter;
  wire             ddr_sdram_clock_crossing_bridge_s1_arb_share_counter_next_value;
  wire             ddr_sdram_clock_crossing_bridge_s1_arb_share_set_values;
  wire             ddr_sdram_clock_crossing_bridge_s1_beginbursttransfer_internal;
  wire             ddr_sdram_clock_crossing_bridge_s1_begins_xfer;
  wire    [  3: 0] ddr_sdram_clock_crossing_bridge_s1_byteenable;
  wire             ddr_sdram_clock_crossing_bridge_s1_end_xfer;
  wire             ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa;
  wire             ddr_sdram_clock_crossing_bridge_s1_firsttransfer;
  wire             ddr_sdram_clock_crossing_bridge_s1_grant_vector;
  wire             ddr_sdram_clock_crossing_bridge_s1_in_a_read_cycle;
  wire             ddr_sdram_clock_crossing_bridge_s1_in_a_write_cycle;
  wire             ddr_sdram_clock_crossing_bridge_s1_master_qreq_vector;
  wire             ddr_sdram_clock_crossing_bridge_s1_move_on_to_next_transaction;
  wire    [ 22: 0] ddr_sdram_clock_crossing_bridge_s1_nativeaddress;
  wire             ddr_sdram_clock_crossing_bridge_s1_non_bursting_master_requests;
  wire             ddr_sdram_clock_crossing_bridge_s1_read;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa;
  wire             ddr_sdram_clock_crossing_bridge_s1_readdatavalid_from_sa;
  reg              ddr_sdram_clock_crossing_bridge_s1_reg_firsttransfer;
  wire             ddr_sdram_clock_crossing_bridge_s1_reset_n;
  reg              ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable;
  wire             ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable2;
  wire             ddr_sdram_clock_crossing_bridge_s1_unreg_firsttransfer;
  wire             ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa;
  wire             ddr_sdram_clock_crossing_bridge_s1_waits_for_read;
  wire             ddr_sdram_clock_crossing_bridge_s1_waits_for_write;
  wire             ddr_sdram_clock_crossing_bridge_s1_write;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_arbiterlock;
  wire             frame_buffer_pipeline_bridge_m1_arbiterlock2;
  wire             frame_buffer_pipeline_bridge_m1_continuerequest;
  wire             frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_rdv_fifo_empty_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_rdv_fifo_output_from_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register;
  wire             frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_saved_grant_ddr_sdram_clock_crossing_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 24: 0] shifted_address_to_ddr_sdram_clock_crossing_bridge_s1_from_frame_buffer_pipeline_bridge_m1;
  wire             wait_for_ddr_sdram_clock_crossing_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ddr_sdram_clock_crossing_bridge_s1_end_xfer;
    end


  assign ddr_sdram_clock_crossing_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1));
  //assign ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa = ddr_sdram_clock_crossing_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa = ddr_sdram_clock_crossing_bridge_s1_readdata;

  assign frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1 = (1) & frame_buffer_pipeline_bridge_m1_chipselect;
  //assign ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa = ddr_sdram_clock_crossing_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa = ddr_sdram_clock_crossing_bridge_s1_waitrequest;

  //assign ddr_sdram_clock_crossing_bridge_s1_readdatavalid_from_sa = ddr_sdram_clock_crossing_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_readdatavalid_from_sa = ddr_sdram_clock_crossing_bridge_s1_readdatavalid;

  //ddr_sdram_clock_crossing_bridge_s1_arb_share_counter set values, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_arb_share_set_values = 1;

  //ddr_sdram_clock_crossing_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_non_bursting_master_requests = frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1;

  //ddr_sdram_clock_crossing_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_any_bursting_master_saved_grant = 0;

  //ddr_sdram_clock_crossing_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_arb_share_counter_next_value = ddr_sdram_clock_crossing_bridge_s1_firsttransfer ? (ddr_sdram_clock_crossing_bridge_s1_arb_share_set_values - 1) : |ddr_sdram_clock_crossing_bridge_s1_arb_share_counter ? (ddr_sdram_clock_crossing_bridge_s1_arb_share_counter - 1) : 0;

  //ddr_sdram_clock_crossing_bridge_s1_allgrants all slave grants, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_allgrants = |ddr_sdram_clock_crossing_bridge_s1_grant_vector;

  //ddr_sdram_clock_crossing_bridge_s1_end_xfer assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_end_xfer = ~(ddr_sdram_clock_crossing_bridge_s1_waits_for_read | ddr_sdram_clock_crossing_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1 = ddr_sdram_clock_crossing_bridge_s1_end_xfer & (~ddr_sdram_clock_crossing_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ddr_sdram_clock_crossing_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1 & ddr_sdram_clock_crossing_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1 & ~ddr_sdram_clock_crossing_bridge_s1_non_bursting_master_requests);

  //ddr_sdram_clock_crossing_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_s1_arb_share_counter <= 0;
      else if (ddr_sdram_clock_crossing_bridge_s1_arb_counter_enable)
          ddr_sdram_clock_crossing_bridge_s1_arb_share_counter <= ddr_sdram_clock_crossing_bridge_s1_arb_share_counter_next_value;
    end


  //ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|ddr_sdram_clock_crossing_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1) | (end_xfer_arb_share_counter_term_ddr_sdram_clock_crossing_bridge_s1 & ~ddr_sdram_clock_crossing_bridge_s1_non_bursting_master_requests))
          ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable <= |ddr_sdram_clock_crossing_bridge_s1_arb_share_counter_next_value;
    end


  //frame_buffer_pipeline_bridge/m1 ddr_sdram_clock_crossing_bridge/s1 arbiterlock, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_arbiterlock = ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable & frame_buffer_pipeline_bridge_m1_continuerequest;

  //ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable2 = |ddr_sdram_clock_crossing_bridge_s1_arb_share_counter_next_value;

  //frame_buffer_pipeline_bridge/m1 ddr_sdram_clock_crossing_bridge/s1 arbiterlock2, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_arbiterlock2 = ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable2 & frame_buffer_pipeline_bridge_m1_continuerequest;

  //ddr_sdram_clock_crossing_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_any_continuerequest = 1;

  //frame_buffer_pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_continuerequest = 1;

  assign frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1 = frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1 & ~(((frame_buffer_pipeline_bridge_m1_read & frame_buffer_pipeline_bridge_m1_chipselect) & ((frame_buffer_pipeline_bridge_m1_latency_counter != 0) | (1 < frame_buffer_pipeline_bridge_m1_latency_counter))));
  //unique name for ddr_sdram_clock_crossing_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_move_on_to_next_transaction = ddr_sdram_clock_crossing_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_frame_buffer_pipeline_bridge_m1_to_ddr_sdram_clock_crossing_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_frame_buffer_pipeline_bridge_m1_to_ddr_sdram_clock_crossing_bridge_s1_module rdv_fifo_for_frame_buffer_pipeline_bridge_m1_to_ddr_sdram_clock_crossing_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1),
      .data_out             (frame_buffer_pipeline_bridge_m1_rdv_fifo_output_from_ddr_sdram_clock_crossing_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (frame_buffer_pipeline_bridge_m1_rdv_fifo_empty_ddr_sdram_clock_crossing_bridge_s1),
      .full                 (),
      .read                 (ddr_sdram_clock_crossing_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr_sdram_clock_crossing_bridge_s1_waits_for_read)
    );

  assign frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register = ~frame_buffer_pipeline_bridge_m1_rdv_fifo_empty_ddr_sdram_clock_crossing_bridge_s1;
  //local readdatavalid frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1, which is an e_mux
  assign frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1 = ddr_sdram_clock_crossing_bridge_s1_readdatavalid_from_sa;

  //ddr_sdram_clock_crossing_bridge_s1_writedata mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_writedata = frame_buffer_pipeline_bridge_m1_writedata;

  //assign ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa = ddr_sdram_clock_crossing_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa = ddr_sdram_clock_crossing_bridge_s1_endofpacket;

  //master is always granted when requested
  assign frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1 = frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1;

  //frame_buffer_pipeline_bridge/m1 saved-grant ddr_sdram_clock_crossing_bridge/s1, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_saved_grant_ddr_sdram_clock_crossing_bridge_s1 = frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1;

  //allow new arb cycle for ddr_sdram_clock_crossing_bridge/s1, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign ddr_sdram_clock_crossing_bridge_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign ddr_sdram_clock_crossing_bridge_s1_master_qreq_vector = 1;

  //ddr_sdram_clock_crossing_bridge_s1_reset_n assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_reset_n = reset_n;

  //ddr_sdram_clock_crossing_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_firsttransfer = ddr_sdram_clock_crossing_bridge_s1_begins_xfer ? ddr_sdram_clock_crossing_bridge_s1_unreg_firsttransfer : ddr_sdram_clock_crossing_bridge_s1_reg_firsttransfer;

  //ddr_sdram_clock_crossing_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_unreg_firsttransfer = ~(ddr_sdram_clock_crossing_bridge_s1_slavearbiterlockenable & ddr_sdram_clock_crossing_bridge_s1_any_continuerequest);

  //ddr_sdram_clock_crossing_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (ddr_sdram_clock_crossing_bridge_s1_begins_xfer)
          ddr_sdram_clock_crossing_bridge_s1_reg_firsttransfer <= ddr_sdram_clock_crossing_bridge_s1_unreg_firsttransfer;
    end


  //ddr_sdram_clock_crossing_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_beginbursttransfer_internal = ddr_sdram_clock_crossing_bridge_s1_begins_xfer;

  //ddr_sdram_clock_crossing_bridge_s1_read assignment, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_read = frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1 & (frame_buffer_pipeline_bridge_m1_read & frame_buffer_pipeline_bridge_m1_chipselect);

  //ddr_sdram_clock_crossing_bridge_s1_write assignment, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_write = frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1 & (frame_buffer_pipeline_bridge_m1_write & frame_buffer_pipeline_bridge_m1_chipselect);

  assign shifted_address_to_ddr_sdram_clock_crossing_bridge_s1_from_frame_buffer_pipeline_bridge_m1 = frame_buffer_pipeline_bridge_m1_address_to_slave;
  //ddr_sdram_clock_crossing_bridge_s1_address mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_address = shifted_address_to_ddr_sdram_clock_crossing_bridge_s1_from_frame_buffer_pipeline_bridge_m1 >> 2;

  //slaveid ddr_sdram_clock_crossing_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_nativeaddress = frame_buffer_pipeline_bridge_m1_address_to_slave >> 2;

  //d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer <= 1;
      else 
        d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer <= ddr_sdram_clock_crossing_bridge_s1_end_xfer;
    end


  //ddr_sdram_clock_crossing_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_waits_for_read = ddr_sdram_clock_crossing_bridge_s1_in_a_read_cycle & ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa;

  //ddr_sdram_clock_crossing_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_in_a_read_cycle = frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1 & (frame_buffer_pipeline_bridge_m1_read & frame_buffer_pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ddr_sdram_clock_crossing_bridge_s1_in_a_read_cycle;

  //ddr_sdram_clock_crossing_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_waits_for_write = ddr_sdram_clock_crossing_bridge_s1_in_a_write_cycle & ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa;

  //ddr_sdram_clock_crossing_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_s1_in_a_write_cycle = frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1 & (frame_buffer_pipeline_bridge_m1_write & frame_buffer_pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ddr_sdram_clock_crossing_bridge_s1_in_a_write_cycle;

  assign wait_for_ddr_sdram_clock_crossing_bridge_s1_counter = 0;
  //ddr_sdram_clock_crossing_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_s1_byteenable = (frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1)? frame_buffer_pipeline_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ddr_sdram_clock_crossing_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //frame_buffer_pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1 && (frame_buffer_pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave ddr_sdram_clock_crossing_bridge/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_clock_crossing_bridge_m1_arbitrator (
                                                       // inputs:
                                                        clk,
                                                        d1_frame_buffer_s1_end_xfer,
                                                        ddr_sdram_clock_crossing_bridge_m1_address,
                                                        ddr_sdram_clock_crossing_bridge_m1_byteenable,
                                                        ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1,
                                                        ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1,
                                                        ddr_sdram_clock_crossing_bridge_m1_read,
                                                        ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1,
                                                        ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register,
                                                        ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1,
                                                        ddr_sdram_clock_crossing_bridge_m1_write,
                                                        ddr_sdram_clock_crossing_bridge_m1_writedata,
                                                        frame_buffer_s1_readdata_from_sa,
                                                        frame_buffer_s1_waitrequest_n_from_sa,
                                                        reset_n,

                                                       // outputs:
                                                        ddr_sdram_clock_crossing_bridge_m1_address_to_slave,
                                                        ddr_sdram_clock_crossing_bridge_m1_latency_counter,
                                                        ddr_sdram_clock_crossing_bridge_m1_readdata,
                                                        ddr_sdram_clock_crossing_bridge_m1_readdatavalid,
                                                        ddr_sdram_clock_crossing_bridge_m1_reset_n,
                                                        ddr_sdram_clock_crossing_bridge_m1_waitrequest
                                                     )
;

  output  [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address_to_slave;
  output           ddr_sdram_clock_crossing_bridge_m1_latency_counter;
  output  [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_readdata;
  output           ddr_sdram_clock_crossing_bridge_m1_readdatavalid;
  output           ddr_sdram_clock_crossing_bridge_m1_reset_n;
  output           ddr_sdram_clock_crossing_bridge_m1_waitrequest;
  input            clk;
  input            d1_frame_buffer_s1_end_xfer;
  input   [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address;
  input   [  3: 0] ddr_sdram_clock_crossing_bridge_m1_byteenable;
  input            ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1;
  input            ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1;
  input            ddr_sdram_clock_crossing_bridge_m1_read;
  input            ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1;
  input            ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register;
  input            ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1;
  input            ddr_sdram_clock_crossing_bridge_m1_write;
  input   [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] frame_buffer_s1_readdata_from_sa;
  input            frame_buffer_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address_last_time;
  wire    [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address_to_slave;
  reg     [  3: 0] ddr_sdram_clock_crossing_bridge_m1_byteenable_last_time;
  wire             ddr_sdram_clock_crossing_bridge_m1_latency_counter;
  reg              ddr_sdram_clock_crossing_bridge_m1_read_last_time;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_readdata;
  wire             ddr_sdram_clock_crossing_bridge_m1_readdatavalid;
  wire             ddr_sdram_clock_crossing_bridge_m1_reset_n;
  wire             ddr_sdram_clock_crossing_bridge_m1_run;
  wire             ddr_sdram_clock_crossing_bridge_m1_waitrequest;
  reg              ddr_sdram_clock_crossing_bridge_m1_write_last_time;
  reg     [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_writedata_last_time;
  wire             pre_flush_ddr_sdram_clock_crossing_bridge_m1_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1 | ~ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1) & ((~ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1 | ~(ddr_sdram_clock_crossing_bridge_m1_read | ddr_sdram_clock_crossing_bridge_m1_write) | (1 & frame_buffer_s1_waitrequest_n_from_sa & (ddr_sdram_clock_crossing_bridge_m1_read | ddr_sdram_clock_crossing_bridge_m1_write)))) & ((~ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1 | ~(ddr_sdram_clock_crossing_bridge_m1_read | ddr_sdram_clock_crossing_bridge_m1_write) | (1 & frame_buffer_s1_waitrequest_n_from_sa & (ddr_sdram_clock_crossing_bridge_m1_read | ddr_sdram_clock_crossing_bridge_m1_write))));

  //cascaded wait assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign ddr_sdram_clock_crossing_bridge_m1_address_to_slave = ddr_sdram_clock_crossing_bridge_m1_address[24 : 0];

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_ddr_sdram_clock_crossing_bridge_m1_readdatavalid = ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_m1_readdatavalid = 0 |
    pre_flush_ddr_sdram_clock_crossing_bridge_m1_readdatavalid;

  //ddr_sdram_clock_crossing_bridge/m1 readdata mux, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_m1_readdata = frame_buffer_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_waitrequest = ~ddr_sdram_clock_crossing_bridge_m1_run;

  //latent max counter, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_latency_counter = 0;

  //ddr_sdram_clock_crossing_bridge_m1_reset_n assignment, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ddr_sdram_clock_crossing_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_m1_address_last_time <= 0;
      else 
        ddr_sdram_clock_crossing_bridge_m1_address_last_time <= ddr_sdram_clock_crossing_bridge_m1_address;
    end


  //ddr_sdram_clock_crossing_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= ddr_sdram_clock_crossing_bridge_m1_waitrequest & (ddr_sdram_clock_crossing_bridge_m1_read | ddr_sdram_clock_crossing_bridge_m1_write);
    end


  //ddr_sdram_clock_crossing_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (ddr_sdram_clock_crossing_bridge_m1_address != ddr_sdram_clock_crossing_bridge_m1_address_last_time))
        begin
          $write("%0d ns: ddr_sdram_clock_crossing_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //ddr_sdram_clock_crossing_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_m1_byteenable_last_time <= 0;
      else 
        ddr_sdram_clock_crossing_bridge_m1_byteenable_last_time <= ddr_sdram_clock_crossing_bridge_m1_byteenable;
    end


  //ddr_sdram_clock_crossing_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (ddr_sdram_clock_crossing_bridge_m1_byteenable != ddr_sdram_clock_crossing_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: ddr_sdram_clock_crossing_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //ddr_sdram_clock_crossing_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_m1_read_last_time <= 0;
      else 
        ddr_sdram_clock_crossing_bridge_m1_read_last_time <= ddr_sdram_clock_crossing_bridge_m1_read;
    end


  //ddr_sdram_clock_crossing_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (ddr_sdram_clock_crossing_bridge_m1_read != ddr_sdram_clock_crossing_bridge_m1_read_last_time))
        begin
          $write("%0d ns: ddr_sdram_clock_crossing_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //ddr_sdram_clock_crossing_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_m1_write_last_time <= 0;
      else 
        ddr_sdram_clock_crossing_bridge_m1_write_last_time <= ddr_sdram_clock_crossing_bridge_m1_write;
    end


  //ddr_sdram_clock_crossing_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (ddr_sdram_clock_crossing_bridge_m1_write != ddr_sdram_clock_crossing_bridge_m1_write_last_time))
        begin
          $write("%0d ns: ddr_sdram_clock_crossing_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //ddr_sdram_clock_crossing_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_clock_crossing_bridge_m1_writedata_last_time <= 0;
      else 
        ddr_sdram_clock_crossing_bridge_m1_writedata_last_time <= ddr_sdram_clock_crossing_bridge_m1_writedata;
    end


  //ddr_sdram_clock_crossing_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (ddr_sdram_clock_crossing_bridge_m1_writedata != ddr_sdram_clock_crossing_bridge_m1_writedata_last_time) & ddr_sdram_clock_crossing_bridge_m1_write)
        begin
          $write("%0d ns: ddr_sdram_clock_crossing_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_clock_crossing_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module descriptor_memory_s1_arbitrator (
                                         // inputs:
                                          clk,
                                          descriptor_memory_s1_readdata,
                                          pipeline_bridge_m1_address_to_slave,
                                          pipeline_bridge_m1_burstcount,
                                          pipeline_bridge_m1_byteenable,
                                          pipeline_bridge_m1_chipselect,
                                          pipeline_bridge_m1_latency_counter,
                                          pipeline_bridge_m1_read,
                                          pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                          pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                          pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                          pipeline_bridge_m1_write,
                                          pipeline_bridge_m1_writedata,
                                          reset_n,

                                         // outputs:
                                          d1_descriptor_memory_s1_end_xfer,
                                          descriptor_memory_s1_address,
                                          descriptor_memory_s1_byteenable,
                                          descriptor_memory_s1_chipselect,
                                          descriptor_memory_s1_clken,
                                          descriptor_memory_s1_readdata_from_sa,
                                          descriptor_memory_s1_reset,
                                          descriptor_memory_s1_write,
                                          descriptor_memory_s1_writedata,
                                          pipeline_bridge_m1_granted_descriptor_memory_s1,
                                          pipeline_bridge_m1_qualified_request_descriptor_memory_s1,
                                          pipeline_bridge_m1_read_data_valid_descriptor_memory_s1,
                                          pipeline_bridge_m1_requests_descriptor_memory_s1
                                       )
;

  output           d1_descriptor_memory_s1_end_xfer;
  output  [  9: 0] descriptor_memory_s1_address;
  output  [  3: 0] descriptor_memory_s1_byteenable;
  output           descriptor_memory_s1_chipselect;
  output           descriptor_memory_s1_clken;
  output  [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  output           descriptor_memory_s1_reset;
  output           descriptor_memory_s1_write;
  output  [ 31: 0] descriptor_memory_s1_writedata;
  output           pipeline_bridge_m1_granted_descriptor_memory_s1;
  output           pipeline_bridge_m1_qualified_request_descriptor_memory_s1;
  output           pipeline_bridge_m1_read_data_valid_descriptor_memory_s1;
  output           pipeline_bridge_m1_requests_descriptor_memory_s1;
  input            clk;
  input   [ 31: 0] descriptor_memory_s1_readdata;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              d1_descriptor_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [  9: 0] descriptor_memory_s1_address;
  wire             descriptor_memory_s1_allgrants;
  wire             descriptor_memory_s1_allow_new_arb_cycle;
  wire             descriptor_memory_s1_any_bursting_master_saved_grant;
  wire             descriptor_memory_s1_any_continuerequest;
  wire             descriptor_memory_s1_arb_counter_enable;
  reg              descriptor_memory_s1_arb_share_counter;
  wire             descriptor_memory_s1_arb_share_counter_next_value;
  wire             descriptor_memory_s1_arb_share_set_values;
  wire             descriptor_memory_s1_beginbursttransfer_internal;
  wire             descriptor_memory_s1_begins_xfer;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire             descriptor_memory_s1_clken;
  wire             descriptor_memory_s1_end_xfer;
  wire             descriptor_memory_s1_firsttransfer;
  wire             descriptor_memory_s1_grant_vector;
  wire             descriptor_memory_s1_in_a_read_cycle;
  wire             descriptor_memory_s1_in_a_write_cycle;
  wire             descriptor_memory_s1_master_qreq_vector;
  wire             descriptor_memory_s1_non_bursting_master_requests;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  reg              descriptor_memory_s1_reg_firsttransfer;
  wire             descriptor_memory_s1_reset;
  reg              descriptor_memory_s1_slavearbiterlockenable;
  wire             descriptor_memory_s1_slavearbiterlockenable2;
  wire             descriptor_memory_s1_unreg_firsttransfer;
  wire             descriptor_memory_s1_waits_for_read;
  wire             descriptor_memory_s1_waits_for_write;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_descriptor_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_descriptor_memory_s1;
  wire             pipeline_bridge_m1_qualified_request_descriptor_memory_s1;
  wire             pipeline_bridge_m1_read_data_valid_descriptor_memory_s1;
  reg              pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register;
  wire             pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             pipeline_bridge_m1_requests_descriptor_memory_s1;
  wire             pipeline_bridge_m1_saved_grant_descriptor_memory_s1;
  wire    [ 26: 0] shifted_address_to_descriptor_memory_s1_from_pipeline_bridge_m1;
  wire             wait_for_descriptor_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~descriptor_memory_s1_end_xfer;
    end


  assign descriptor_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_descriptor_memory_s1));
  //assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata;

  assign pipeline_bridge_m1_requests_descriptor_memory_s1 = ({pipeline_bridge_m1_address_to_slave[26 : 12] , 12'b0} == 27'h4400000) & pipeline_bridge_m1_chipselect;
  //descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  assign descriptor_memory_s1_arb_share_set_values = 1;

  //descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign descriptor_memory_s1_non_bursting_master_requests = pipeline_bridge_m1_requests_descriptor_memory_s1;

  //descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign descriptor_memory_s1_any_bursting_master_saved_grant = 0;

  //descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign descriptor_memory_s1_arb_share_counter_next_value = descriptor_memory_s1_firsttransfer ? (descriptor_memory_s1_arb_share_set_values - 1) : |descriptor_memory_s1_arb_share_counter ? (descriptor_memory_s1_arb_share_counter - 1) : 0;

  //descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  assign descriptor_memory_s1_allgrants = |descriptor_memory_s1_grant_vector;

  //descriptor_memory_s1_end_xfer assignment, which is an e_assign
  assign descriptor_memory_s1_end_xfer = ~(descriptor_memory_s1_waits_for_read | descriptor_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_descriptor_memory_s1 = descriptor_memory_s1_end_xfer & (~descriptor_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign descriptor_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_descriptor_memory_s1 & descriptor_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests);

  //descriptor_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_share_counter <= 0;
      else if (descriptor_memory_s1_arb_counter_enable)
          descriptor_memory_s1_arb_share_counter <= descriptor_memory_s1_arb_share_counter_next_value;
    end


  //descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_slavearbiterlockenable <= 0;
      else if ((|descriptor_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_descriptor_memory_s1) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests))
          descriptor_memory_s1_slavearbiterlockenable <= |descriptor_memory_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 descriptor_memory/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign descriptor_memory_s1_slavearbiterlockenable2 = |descriptor_memory_s1_arb_share_counter_next_value;

  //pipeline_bridge/m1 descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign descriptor_memory_s1_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_descriptor_memory_s1 = pipeline_bridge_m1_requests_descriptor_memory_s1 & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((1 < pipeline_bridge_m1_latency_counter) | (|pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register))));
  //pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in = pipeline_bridge_m1_granted_descriptor_memory_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register = {pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register, pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in};

  //pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register <= p1_pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid pipeline_bridge_m1_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_descriptor_memory_s1 = pipeline_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register;

  //descriptor_memory_s1_writedata mux, which is an e_mux
  assign descriptor_memory_s1_writedata = pipeline_bridge_m1_writedata;

  //mux descriptor_memory_s1_clken, which is an e_mux
  assign descriptor_memory_s1_clken = 1'b1;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_descriptor_memory_s1 = pipeline_bridge_m1_qualified_request_descriptor_memory_s1;

  //pipeline_bridge/m1 saved-grant descriptor_memory/s1, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_descriptor_memory_s1 = pipeline_bridge_m1_requests_descriptor_memory_s1;

  //allow new arb cycle for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign descriptor_memory_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign descriptor_memory_s1_master_qreq_vector = 1;

  //~descriptor_memory_s1_reset assignment, which is an e_assign
  assign descriptor_memory_s1_reset = ~reset_n;

  assign descriptor_memory_s1_chipselect = pipeline_bridge_m1_granted_descriptor_memory_s1;
  //descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_firsttransfer = descriptor_memory_s1_begins_xfer ? descriptor_memory_s1_unreg_firsttransfer : descriptor_memory_s1_reg_firsttransfer;

  //descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_unreg_firsttransfer = ~(descriptor_memory_s1_slavearbiterlockenable & descriptor_memory_s1_any_continuerequest);

  //descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_reg_firsttransfer <= 1'b1;
      else if (descriptor_memory_s1_begins_xfer)
          descriptor_memory_s1_reg_firsttransfer <= descriptor_memory_s1_unreg_firsttransfer;
    end


  //descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign descriptor_memory_s1_beginbursttransfer_internal = descriptor_memory_s1_begins_xfer;

  //descriptor_memory_s1_write assignment, which is an e_mux
  assign descriptor_memory_s1_write = pipeline_bridge_m1_granted_descriptor_memory_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_descriptor_memory_s1_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //descriptor_memory_s1_address mux, which is an e_mux
  assign descriptor_memory_s1_address = shifted_address_to_descriptor_memory_s1_from_pipeline_bridge_m1 >> 2;

  //d1_descriptor_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_descriptor_memory_s1_end_xfer <= 1;
      else 
        d1_descriptor_memory_s1_end_xfer <= descriptor_memory_s1_end_xfer;
    end


  //descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_read = descriptor_memory_s1_in_a_read_cycle & 0;

  //descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_read_cycle = pipeline_bridge_m1_granted_descriptor_memory_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = descriptor_memory_s1_in_a_read_cycle;

  //descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_write = descriptor_memory_s1_in_a_write_cycle & 0;

  //descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_write_cycle = pipeline_bridge_m1_granted_descriptor_memory_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = descriptor_memory_s1_in_a_write_cycle;

  assign wait_for_descriptor_memory_s1_counter = 0;
  //descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign descriptor_memory_s1_byteenable = (pipeline_bridge_m1_granted_descriptor_memory_s1)? pipeline_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //descriptor_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_descriptor_memory_s1 && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave descriptor_memory/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module descriptor_memory_s2_arbitrator (
                                         // inputs:
                                          clk,
                                          descriptor_memory_s2_readdata,
                                          lcd_sgdma_descriptor_read_address_to_slave,
                                          lcd_sgdma_descriptor_read_latency_counter,
                                          lcd_sgdma_descriptor_read_read,
                                          lcd_sgdma_descriptor_write_address_to_slave,
                                          lcd_sgdma_descriptor_write_write,
                                          lcd_sgdma_descriptor_write_writedata,
                                          reset_n,

                                         // outputs:
                                          d1_descriptor_memory_s2_end_xfer,
                                          descriptor_memory_s2_address,
                                          descriptor_memory_s2_byteenable,
                                          descriptor_memory_s2_chipselect,
                                          descriptor_memory_s2_clken,
                                          descriptor_memory_s2_readdata_from_sa,
                                          descriptor_memory_s2_reset,
                                          descriptor_memory_s2_write,
                                          descriptor_memory_s2_writedata,
                                          lcd_sgdma_descriptor_read_granted_descriptor_memory_s2,
                                          lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2,
                                          lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2,
                                          lcd_sgdma_descriptor_read_requests_descriptor_memory_s2,
                                          lcd_sgdma_descriptor_write_granted_descriptor_memory_s2,
                                          lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2,
                                          lcd_sgdma_descriptor_write_requests_descriptor_memory_s2
                                       )
;

  output           d1_descriptor_memory_s2_end_xfer;
  output  [  9: 0] descriptor_memory_s2_address;
  output  [  3: 0] descriptor_memory_s2_byteenable;
  output           descriptor_memory_s2_chipselect;
  output           descriptor_memory_s2_clken;
  output  [ 31: 0] descriptor_memory_s2_readdata_from_sa;
  output           descriptor_memory_s2_reset;
  output           descriptor_memory_s2_write;
  output  [ 31: 0] descriptor_memory_s2_writedata;
  output           lcd_sgdma_descriptor_read_granted_descriptor_memory_s2;
  output           lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2;
  output           lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2;
  output           lcd_sgdma_descriptor_read_requests_descriptor_memory_s2;
  output           lcd_sgdma_descriptor_write_granted_descriptor_memory_s2;
  output           lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2;
  output           lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;
  input            clk;
  input   [ 31: 0] descriptor_memory_s2_readdata;
  input   [ 31: 0] lcd_sgdma_descriptor_read_address_to_slave;
  input            lcd_sgdma_descriptor_read_latency_counter;
  input            lcd_sgdma_descriptor_read_read;
  input   [ 31: 0] lcd_sgdma_descriptor_write_address_to_slave;
  input            lcd_sgdma_descriptor_write_write;
  input   [ 31: 0] lcd_sgdma_descriptor_write_writedata;
  input            reset_n;

  reg              d1_descriptor_memory_s2_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [  9: 0] descriptor_memory_s2_address;
  wire             descriptor_memory_s2_allgrants;
  wire             descriptor_memory_s2_allow_new_arb_cycle;
  wire             descriptor_memory_s2_any_bursting_master_saved_grant;
  wire             descriptor_memory_s2_any_continuerequest;
  reg     [  1: 0] descriptor_memory_s2_arb_addend;
  wire             descriptor_memory_s2_arb_counter_enable;
  reg              descriptor_memory_s2_arb_share_counter;
  wire             descriptor_memory_s2_arb_share_counter_next_value;
  wire             descriptor_memory_s2_arb_share_set_values;
  wire    [  1: 0] descriptor_memory_s2_arb_winner;
  wire             descriptor_memory_s2_arbitration_holdoff_internal;
  wire             descriptor_memory_s2_beginbursttransfer_internal;
  wire             descriptor_memory_s2_begins_xfer;
  wire    [  3: 0] descriptor_memory_s2_byteenable;
  wire             descriptor_memory_s2_chipselect;
  wire    [  3: 0] descriptor_memory_s2_chosen_master_double_vector;
  wire    [  1: 0] descriptor_memory_s2_chosen_master_rot_left;
  wire             descriptor_memory_s2_clken;
  wire             descriptor_memory_s2_end_xfer;
  wire             descriptor_memory_s2_firsttransfer;
  wire    [  1: 0] descriptor_memory_s2_grant_vector;
  wire             descriptor_memory_s2_in_a_read_cycle;
  wire             descriptor_memory_s2_in_a_write_cycle;
  wire    [  1: 0] descriptor_memory_s2_master_qreq_vector;
  wire             descriptor_memory_s2_non_bursting_master_requests;
  wire    [ 31: 0] descriptor_memory_s2_readdata_from_sa;
  reg              descriptor_memory_s2_reg_firsttransfer;
  wire             descriptor_memory_s2_reset;
  reg     [  1: 0] descriptor_memory_s2_saved_chosen_master_vector;
  reg              descriptor_memory_s2_slavearbiterlockenable;
  wire             descriptor_memory_s2_slavearbiterlockenable2;
  wire             descriptor_memory_s2_unreg_firsttransfer;
  wire             descriptor_memory_s2_waits_for_read;
  wire             descriptor_memory_s2_waits_for_write;
  wire             descriptor_memory_s2_write;
  wire    [ 31: 0] descriptor_memory_s2_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_descriptor_memory_s2;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_lcd_sgdma_descriptor_read_granted_slave_descriptor_memory_s2;
  reg              last_cycle_lcd_sgdma_descriptor_write_granted_slave_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_arbiterlock;
  wire             lcd_sgdma_descriptor_read_arbiterlock2;
  wire             lcd_sgdma_descriptor_read_continuerequest;
  wire             lcd_sgdma_descriptor_read_granted_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2;
  reg              lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register;
  wire             lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register_in;
  wire             lcd_sgdma_descriptor_read_requests_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_saved_grant_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_arbiterlock;
  wire             lcd_sgdma_descriptor_write_arbiterlock2;
  wire             lcd_sgdma_descriptor_write_continuerequest;
  wire             lcd_sgdma_descriptor_write_granted_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_saved_grant_descriptor_memory_s2;
  wire             p1_lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s2_from_lcd_sgdma_descriptor_read;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s2_from_lcd_sgdma_descriptor_write;
  wire             wait_for_descriptor_memory_s2_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~descriptor_memory_s2_end_xfer;
    end


  assign descriptor_memory_s2_begins_xfer = ~d1_reasons_to_wait & ((lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2 | lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2));
  //assign descriptor_memory_s2_readdata_from_sa = descriptor_memory_s2_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign descriptor_memory_s2_readdata_from_sa = descriptor_memory_s2_readdata;

  assign lcd_sgdma_descriptor_read_requests_descriptor_memory_s2 = (({lcd_sgdma_descriptor_read_address_to_slave[31 : 12] , 12'b0} == 32'h4400000) & (lcd_sgdma_descriptor_read_read)) & lcd_sgdma_descriptor_read_read;
  //descriptor_memory_s2_arb_share_counter set values, which is an e_mux
  assign descriptor_memory_s2_arb_share_set_values = 1;

  //descriptor_memory_s2_non_bursting_master_requests mux, which is an e_mux
  assign descriptor_memory_s2_non_bursting_master_requests = lcd_sgdma_descriptor_read_requests_descriptor_memory_s2 |
    lcd_sgdma_descriptor_write_requests_descriptor_memory_s2 |
    lcd_sgdma_descriptor_read_requests_descriptor_memory_s2 |
    lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;

  //descriptor_memory_s2_any_bursting_master_saved_grant mux, which is an e_mux
  assign descriptor_memory_s2_any_bursting_master_saved_grant = 0;

  //descriptor_memory_s2_arb_share_counter_next_value assignment, which is an e_assign
  assign descriptor_memory_s2_arb_share_counter_next_value = descriptor_memory_s2_firsttransfer ? (descriptor_memory_s2_arb_share_set_values - 1) : |descriptor_memory_s2_arb_share_counter ? (descriptor_memory_s2_arb_share_counter - 1) : 0;

  //descriptor_memory_s2_allgrants all slave grants, which is an e_mux
  assign descriptor_memory_s2_allgrants = (|descriptor_memory_s2_grant_vector) |
    (|descriptor_memory_s2_grant_vector) |
    (|descriptor_memory_s2_grant_vector) |
    (|descriptor_memory_s2_grant_vector);

  //descriptor_memory_s2_end_xfer assignment, which is an e_assign
  assign descriptor_memory_s2_end_xfer = ~(descriptor_memory_s2_waits_for_read | descriptor_memory_s2_waits_for_write);

  //end_xfer_arb_share_counter_term_descriptor_memory_s2 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_descriptor_memory_s2 = descriptor_memory_s2_end_xfer & (~descriptor_memory_s2_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //descriptor_memory_s2_arb_share_counter arbitration counter enable, which is an e_assign
  assign descriptor_memory_s2_arb_counter_enable = (end_xfer_arb_share_counter_term_descriptor_memory_s2 & descriptor_memory_s2_allgrants) | (end_xfer_arb_share_counter_term_descriptor_memory_s2 & ~descriptor_memory_s2_non_bursting_master_requests);

  //descriptor_memory_s2_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s2_arb_share_counter <= 0;
      else if (descriptor_memory_s2_arb_counter_enable)
          descriptor_memory_s2_arb_share_counter <= descriptor_memory_s2_arb_share_counter_next_value;
    end


  //descriptor_memory_s2_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s2_slavearbiterlockenable <= 0;
      else if ((|descriptor_memory_s2_master_qreq_vector & end_xfer_arb_share_counter_term_descriptor_memory_s2) | (end_xfer_arb_share_counter_term_descriptor_memory_s2 & ~descriptor_memory_s2_non_bursting_master_requests))
          descriptor_memory_s2_slavearbiterlockenable <= |descriptor_memory_s2_arb_share_counter_next_value;
    end


  //lcd_sgdma/descriptor_read descriptor_memory/s2 arbiterlock, which is an e_assign
  assign lcd_sgdma_descriptor_read_arbiterlock = descriptor_memory_s2_slavearbiterlockenable & lcd_sgdma_descriptor_read_continuerequest;

  //descriptor_memory_s2_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign descriptor_memory_s2_slavearbiterlockenable2 = |descriptor_memory_s2_arb_share_counter_next_value;

  //lcd_sgdma/descriptor_read descriptor_memory/s2 arbiterlock2, which is an e_assign
  assign lcd_sgdma_descriptor_read_arbiterlock2 = descriptor_memory_s2_slavearbiterlockenable2 & lcd_sgdma_descriptor_read_continuerequest;

  //lcd_sgdma/descriptor_write descriptor_memory/s2 arbiterlock, which is an e_assign
  assign lcd_sgdma_descriptor_write_arbiterlock = descriptor_memory_s2_slavearbiterlockenable & lcd_sgdma_descriptor_write_continuerequest;

  //lcd_sgdma/descriptor_write descriptor_memory/s2 arbiterlock2, which is an e_assign
  assign lcd_sgdma_descriptor_write_arbiterlock2 = descriptor_memory_s2_slavearbiterlockenable2 & lcd_sgdma_descriptor_write_continuerequest;

  //lcd_sgdma/descriptor_write granted descriptor_memory/s2 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_lcd_sgdma_descriptor_write_granted_slave_descriptor_memory_s2 <= 0;
      else 
        last_cycle_lcd_sgdma_descriptor_write_granted_slave_descriptor_memory_s2 <= lcd_sgdma_descriptor_write_saved_grant_descriptor_memory_s2 ? 1 : (descriptor_memory_s2_arbitration_holdoff_internal | ~lcd_sgdma_descriptor_write_requests_descriptor_memory_s2) ? 0 : last_cycle_lcd_sgdma_descriptor_write_granted_slave_descriptor_memory_s2;
    end


  //lcd_sgdma_descriptor_write_continuerequest continued request, which is an e_mux
  assign lcd_sgdma_descriptor_write_continuerequest = last_cycle_lcd_sgdma_descriptor_write_granted_slave_descriptor_memory_s2 & lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;

  //descriptor_memory_s2_any_continuerequest at least one master continues requesting, which is an e_mux
  assign descriptor_memory_s2_any_continuerequest = lcd_sgdma_descriptor_write_continuerequest |
    lcd_sgdma_descriptor_read_continuerequest;

  assign lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2 = lcd_sgdma_descriptor_read_requests_descriptor_memory_s2 & ~(lcd_sgdma_descriptor_write_arbiterlock);
  //lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register_in mux for readlatency shift register, which is an e_mux
  assign lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register_in = lcd_sgdma_descriptor_read_granted_descriptor_memory_s2 & lcd_sgdma_descriptor_read_read & ~descriptor_memory_s2_waits_for_read;

  //shift register p1 lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register = {lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register, lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register_in};

  //lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register <= 0;
      else 
        lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register <= p1_lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register;
    end


  //local readdatavalid lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2, which is an e_mux
  assign lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2 = lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2_shift_register;

  //mux descriptor_memory_s2_clken, which is an e_mux
  assign descriptor_memory_s2_clken = 1'b1;

  assign lcd_sgdma_descriptor_write_requests_descriptor_memory_s2 = (({lcd_sgdma_descriptor_write_address_to_slave[31 : 12] , 12'b0} == 32'h4400000) & (lcd_sgdma_descriptor_write_write)) & lcd_sgdma_descriptor_write_write;
  //lcd_sgdma/descriptor_read granted descriptor_memory/s2 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_lcd_sgdma_descriptor_read_granted_slave_descriptor_memory_s2 <= 0;
      else 
        last_cycle_lcd_sgdma_descriptor_read_granted_slave_descriptor_memory_s2 <= lcd_sgdma_descriptor_read_saved_grant_descriptor_memory_s2 ? 1 : (descriptor_memory_s2_arbitration_holdoff_internal | ~lcd_sgdma_descriptor_read_requests_descriptor_memory_s2) ? 0 : last_cycle_lcd_sgdma_descriptor_read_granted_slave_descriptor_memory_s2;
    end


  //lcd_sgdma_descriptor_read_continuerequest continued request, which is an e_mux
  assign lcd_sgdma_descriptor_read_continuerequest = last_cycle_lcd_sgdma_descriptor_read_granted_slave_descriptor_memory_s2 & lcd_sgdma_descriptor_read_requests_descriptor_memory_s2;

  assign lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2 = lcd_sgdma_descriptor_write_requests_descriptor_memory_s2 & ~(lcd_sgdma_descriptor_read_arbiterlock);
  //descriptor_memory_s2_writedata mux, which is an e_mux
  assign descriptor_memory_s2_writedata = lcd_sgdma_descriptor_write_writedata;

  //allow new arb cycle for descriptor_memory/s2, which is an e_assign
  assign descriptor_memory_s2_allow_new_arb_cycle = ~lcd_sgdma_descriptor_read_arbiterlock & ~lcd_sgdma_descriptor_write_arbiterlock;

  //lcd_sgdma/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s2, which is an e_assign
  assign descriptor_memory_s2_master_qreq_vector[0] = lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2;

  //lcd_sgdma/descriptor_write grant descriptor_memory/s2, which is an e_assign
  assign lcd_sgdma_descriptor_write_granted_descriptor_memory_s2 = descriptor_memory_s2_grant_vector[0];

  //lcd_sgdma/descriptor_write saved-grant descriptor_memory/s2, which is an e_assign
  assign lcd_sgdma_descriptor_write_saved_grant_descriptor_memory_s2 = descriptor_memory_s2_arb_winner[0] && lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;

  //lcd_sgdma/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s2, which is an e_assign
  assign descriptor_memory_s2_master_qreq_vector[1] = lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2;

  //lcd_sgdma/descriptor_read grant descriptor_memory/s2, which is an e_assign
  assign lcd_sgdma_descriptor_read_granted_descriptor_memory_s2 = descriptor_memory_s2_grant_vector[1];

  //lcd_sgdma/descriptor_read saved-grant descriptor_memory/s2, which is an e_assign
  assign lcd_sgdma_descriptor_read_saved_grant_descriptor_memory_s2 = descriptor_memory_s2_arb_winner[1] && lcd_sgdma_descriptor_read_requests_descriptor_memory_s2;

  //descriptor_memory/s2 chosen-master double-vector, which is an e_assign
  assign descriptor_memory_s2_chosen_master_double_vector = {descriptor_memory_s2_master_qreq_vector, descriptor_memory_s2_master_qreq_vector} & ({~descriptor_memory_s2_master_qreq_vector, ~descriptor_memory_s2_master_qreq_vector} + descriptor_memory_s2_arb_addend);

  //stable onehot encoding of arb winner
  assign descriptor_memory_s2_arb_winner = (descriptor_memory_s2_allow_new_arb_cycle & | descriptor_memory_s2_grant_vector) ? descriptor_memory_s2_grant_vector : descriptor_memory_s2_saved_chosen_master_vector;

  //saved descriptor_memory_s2_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s2_saved_chosen_master_vector <= 0;
      else if (descriptor_memory_s2_allow_new_arb_cycle)
          descriptor_memory_s2_saved_chosen_master_vector <= |descriptor_memory_s2_grant_vector ? descriptor_memory_s2_grant_vector : descriptor_memory_s2_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign descriptor_memory_s2_grant_vector = {(descriptor_memory_s2_chosen_master_double_vector[1] | descriptor_memory_s2_chosen_master_double_vector[3]),
    (descriptor_memory_s2_chosen_master_double_vector[0] | descriptor_memory_s2_chosen_master_double_vector[2])};

  //descriptor_memory/s2 chosen master rotated left, which is an e_assign
  assign descriptor_memory_s2_chosen_master_rot_left = (descriptor_memory_s2_arb_winner << 1) ? (descriptor_memory_s2_arb_winner << 1) : 1;

  //descriptor_memory/s2's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s2_arb_addend <= 1;
      else if (|descriptor_memory_s2_grant_vector)
          descriptor_memory_s2_arb_addend <= descriptor_memory_s2_end_xfer? descriptor_memory_s2_chosen_master_rot_left : descriptor_memory_s2_grant_vector;
    end


  //~descriptor_memory_s2_reset assignment, which is an e_assign
  assign descriptor_memory_s2_reset = ~reset_n;

  assign descriptor_memory_s2_chipselect = lcd_sgdma_descriptor_read_granted_descriptor_memory_s2 | lcd_sgdma_descriptor_write_granted_descriptor_memory_s2;
  //descriptor_memory_s2_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s2_firsttransfer = descriptor_memory_s2_begins_xfer ? descriptor_memory_s2_unreg_firsttransfer : descriptor_memory_s2_reg_firsttransfer;

  //descriptor_memory_s2_unreg_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s2_unreg_firsttransfer = ~(descriptor_memory_s2_slavearbiterlockenable & descriptor_memory_s2_any_continuerequest);

  //descriptor_memory_s2_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s2_reg_firsttransfer <= 1'b1;
      else if (descriptor_memory_s2_begins_xfer)
          descriptor_memory_s2_reg_firsttransfer <= descriptor_memory_s2_unreg_firsttransfer;
    end


  //descriptor_memory_s2_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign descriptor_memory_s2_beginbursttransfer_internal = descriptor_memory_s2_begins_xfer;

  //descriptor_memory_s2_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign descriptor_memory_s2_arbitration_holdoff_internal = descriptor_memory_s2_begins_xfer & descriptor_memory_s2_firsttransfer;

  //descriptor_memory_s2_write assignment, which is an e_mux
  assign descriptor_memory_s2_write = lcd_sgdma_descriptor_write_granted_descriptor_memory_s2 & lcd_sgdma_descriptor_write_write;

  assign shifted_address_to_descriptor_memory_s2_from_lcd_sgdma_descriptor_read = lcd_sgdma_descriptor_read_address_to_slave;
  //descriptor_memory_s2_address mux, which is an e_mux
  assign descriptor_memory_s2_address = (lcd_sgdma_descriptor_read_granted_descriptor_memory_s2)? (shifted_address_to_descriptor_memory_s2_from_lcd_sgdma_descriptor_read >> 2) :
    (shifted_address_to_descriptor_memory_s2_from_lcd_sgdma_descriptor_write >> 2);

  assign shifted_address_to_descriptor_memory_s2_from_lcd_sgdma_descriptor_write = lcd_sgdma_descriptor_write_address_to_slave;
  //d1_descriptor_memory_s2_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_descriptor_memory_s2_end_xfer <= 1;
      else 
        d1_descriptor_memory_s2_end_xfer <= descriptor_memory_s2_end_xfer;
    end


  //descriptor_memory_s2_waits_for_read in a cycle, which is an e_mux
  assign descriptor_memory_s2_waits_for_read = descriptor_memory_s2_in_a_read_cycle & 0;

  //descriptor_memory_s2_in_a_read_cycle assignment, which is an e_assign
  assign descriptor_memory_s2_in_a_read_cycle = lcd_sgdma_descriptor_read_granted_descriptor_memory_s2 & lcd_sgdma_descriptor_read_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = descriptor_memory_s2_in_a_read_cycle;

  //descriptor_memory_s2_waits_for_write in a cycle, which is an e_mux
  assign descriptor_memory_s2_waits_for_write = descriptor_memory_s2_in_a_write_cycle & 0;

  //descriptor_memory_s2_in_a_write_cycle assignment, which is an e_assign
  assign descriptor_memory_s2_in_a_write_cycle = lcd_sgdma_descriptor_write_granted_descriptor_memory_s2 & lcd_sgdma_descriptor_write_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = descriptor_memory_s2_in_a_write_cycle;

  assign wait_for_descriptor_memory_s2_counter = 0;
  //descriptor_memory_s2_byteenable byte enable port mux, which is an e_mux
  assign descriptor_memory_s2_byteenable = (lcd_sgdma_descriptor_write_granted_descriptor_memory_s2)? {4 {1'b1}} :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //descriptor_memory/s2 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (lcd_sgdma_descriptor_read_granted_descriptor_memory_s2 + lcd_sgdma_descriptor_write_granted_descriptor_memory_s2 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (lcd_sgdma_descriptor_read_saved_grant_descriptor_memory_s2 + lcd_sgdma_descriptor_write_saved_grant_descriptor_memory_s2 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module dummy_master_inst_m0_arbitrator (
                                         // inputs:
                                          clk,
                                          d1_colour_lookup_table_s2_end_xfer,
                                          dummy_master_inst_granted_colour_lookup_table_s2,
                                          dummy_master_inst_m0_address,
                                          dummy_master_inst_m0_write,
                                          dummy_master_inst_m0_writedata,
                                          dummy_master_inst_qualified_request_colour_lookup_table_s2,
                                          dummy_master_inst_requests_colour_lookup_table_s2,
                                          reset_n,

                                         // outputs:
                                          dummy_master_inst_m0_address_to_slave,
                                          dummy_master_inst_m0_waitrequest
                                       )
;

  output  [ 31: 0] dummy_master_inst_m0_address_to_slave;
  output           dummy_master_inst_m0_waitrequest;
  input            clk;
  input            d1_colour_lookup_table_s2_end_xfer;
  input            dummy_master_inst_granted_colour_lookup_table_s2;
  input   [ 31: 0] dummy_master_inst_m0_address;
  input            dummy_master_inst_m0_write;
  input   [ 31: 0] dummy_master_inst_m0_writedata;
  input            dummy_master_inst_qualified_request_colour_lookup_table_s2;
  input            dummy_master_inst_requests_colour_lookup_table_s2;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 31: 0] dummy_master_inst_m0_address_last_time;
  wire    [ 31: 0] dummy_master_inst_m0_address_to_slave;
  wire             dummy_master_inst_m0_run;
  wire             dummy_master_inst_m0_waitrequest;
  reg              dummy_master_inst_m0_write_last_time;
  reg     [ 31: 0] dummy_master_inst_m0_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (dummy_master_inst_qualified_request_colour_lookup_table_s2 | ~dummy_master_inst_requests_colour_lookup_table_s2) & (dummy_master_inst_granted_colour_lookup_table_s2 | ~dummy_master_inst_qualified_request_colour_lookup_table_s2) & ((~dummy_master_inst_qualified_request_colour_lookup_table_s2 | ~(dummy_master_inst_m0_write) | (1 & (dummy_master_inst_m0_write))));

  //cascaded wait assignment, which is an e_assign
  assign dummy_master_inst_m0_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign dummy_master_inst_m0_address_to_slave = {22'b10001000000000111,
    dummy_master_inst_m0_address[9 : 0]};

  //actual waitrequest port, which is an e_assign
  assign dummy_master_inst_m0_waitrequest = ~dummy_master_inst_m0_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //dummy_master_inst_m0_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dummy_master_inst_m0_address_last_time <= 0;
      else 
        dummy_master_inst_m0_address_last_time <= dummy_master_inst_m0_address;
    end


  //dummy_master_inst/m0 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= dummy_master_inst_m0_waitrequest & (dummy_master_inst_m0_write);
    end


  //dummy_master_inst_m0_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (dummy_master_inst_m0_address != dummy_master_inst_m0_address_last_time))
        begin
          $write("%0d ns: dummy_master_inst_m0_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //dummy_master_inst_m0_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dummy_master_inst_m0_write_last_time <= 0;
      else 
        dummy_master_inst_m0_write_last_time <= dummy_master_inst_m0_write;
    end


  //dummy_master_inst_m0_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (dummy_master_inst_m0_write != dummy_master_inst_m0_write_last_time))
        begin
          $write("%0d ns: dummy_master_inst_m0_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //dummy_master_inst_m0_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dummy_master_inst_m0_writedata_last_time <= 0;
      else 
        dummy_master_inst_m0_writedata_last_time <= dummy_master_inst_m0_writedata;
    end


  //dummy_master_inst_m0_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (dummy_master_inst_m0_writedata != dummy_master_inst_m0_writedata_last_time) & dummy_master_inst_m0_write)
        begin
          $write("%0d ns: dummy_master_inst_m0_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_pipeline_bridge_m1_to_flash_ssram_pipeline_bridge_s1_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_ssram_pipeline_bridge_s1_arbitrator (
                                                   // inputs:
                                                    clk,
                                                    flash_ssram_pipeline_bridge_s1_endofpacket,
                                                    flash_ssram_pipeline_bridge_s1_readdata,
                                                    flash_ssram_pipeline_bridge_s1_readdatavalid,
                                                    flash_ssram_pipeline_bridge_s1_waitrequest,
                                                    pipeline_bridge_m1_address_to_slave,
                                                    pipeline_bridge_m1_burstcount,
                                                    pipeline_bridge_m1_byteenable,
                                                    pipeline_bridge_m1_chipselect,
                                                    pipeline_bridge_m1_debugaccess,
                                                    pipeline_bridge_m1_latency_counter,
                                                    pipeline_bridge_m1_read,
                                                    pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                                    pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                                    pipeline_bridge_m1_write,
                                                    pipeline_bridge_m1_writedata,
                                                    reset_n,

                                                   // outputs:
                                                    d1_flash_ssram_pipeline_bridge_s1_end_xfer,
                                                    flash_ssram_pipeline_bridge_s1_address,
                                                    flash_ssram_pipeline_bridge_s1_arbiterlock,
                                                    flash_ssram_pipeline_bridge_s1_arbiterlock2,
                                                    flash_ssram_pipeline_bridge_s1_burstcount,
                                                    flash_ssram_pipeline_bridge_s1_byteenable,
                                                    flash_ssram_pipeline_bridge_s1_chipselect,
                                                    flash_ssram_pipeline_bridge_s1_debugaccess,
                                                    flash_ssram_pipeline_bridge_s1_endofpacket_from_sa,
                                                    flash_ssram_pipeline_bridge_s1_nativeaddress,
                                                    flash_ssram_pipeline_bridge_s1_read,
                                                    flash_ssram_pipeline_bridge_s1_readdata_from_sa,
                                                    flash_ssram_pipeline_bridge_s1_reset_n,
                                                    flash_ssram_pipeline_bridge_s1_waitrequest_from_sa,
                                                    flash_ssram_pipeline_bridge_s1_write,
                                                    flash_ssram_pipeline_bridge_s1_writedata,
                                                    pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1,
                                                    pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1,
                                                    pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1,
                                                    pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                                    pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1
                                                 )
;

  output           d1_flash_ssram_pipeline_bridge_s1_end_xfer;
  output  [ 19: 0] flash_ssram_pipeline_bridge_s1_address;
  output           flash_ssram_pipeline_bridge_s1_arbiterlock;
  output           flash_ssram_pipeline_bridge_s1_arbiterlock2;
  output           flash_ssram_pipeline_bridge_s1_burstcount;
  output  [ 31: 0] flash_ssram_pipeline_bridge_s1_byteenable;
  output           flash_ssram_pipeline_bridge_s1_chipselect;
  output           flash_ssram_pipeline_bridge_s1_debugaccess;
  output           flash_ssram_pipeline_bridge_s1_endofpacket_from_sa;
  output  [ 19: 0] flash_ssram_pipeline_bridge_s1_nativeaddress;
  output           flash_ssram_pipeline_bridge_s1_read;
  output  [255: 0] flash_ssram_pipeline_bridge_s1_readdata_from_sa;
  output           flash_ssram_pipeline_bridge_s1_reset_n;
  output           flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
  output           flash_ssram_pipeline_bridge_s1_write;
  output  [255: 0] flash_ssram_pipeline_bridge_s1_writedata;
  output           pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1;
  output           pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1;
  output           pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1;
  output           pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  output           pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;
  input            clk;
  input            flash_ssram_pipeline_bridge_s1_endofpacket;
  input   [255: 0] flash_ssram_pipeline_bridge_s1_readdata;
  input            flash_ssram_pipeline_bridge_s1_readdatavalid;
  input            flash_ssram_pipeline_bridge_s1_waitrequest;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_debugaccess;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              d1_flash_ssram_pipeline_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1;
  wire    [ 19: 0] flash_ssram_pipeline_bridge_s1_address;
  wire             flash_ssram_pipeline_bridge_s1_allgrants;
  wire             flash_ssram_pipeline_bridge_s1_allow_new_arb_cycle;
  wire             flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant;
  wire             flash_ssram_pipeline_bridge_s1_any_continuerequest;
  wire             flash_ssram_pipeline_bridge_s1_arb_counter_enable;
  reg              flash_ssram_pipeline_bridge_s1_arb_share_counter;
  wire             flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;
  wire             flash_ssram_pipeline_bridge_s1_arb_share_set_values;
  wire             flash_ssram_pipeline_bridge_s1_arbiterlock;
  wire             flash_ssram_pipeline_bridge_s1_arbiterlock2;
  wire             flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal;
  wire             flash_ssram_pipeline_bridge_s1_beginbursttransfer_internal;
  wire             flash_ssram_pipeline_bridge_s1_begins_xfer;
  wire             flash_ssram_pipeline_bridge_s1_burstcount;
  wire    [ 31: 0] flash_ssram_pipeline_bridge_s1_byteenable;
  wire             flash_ssram_pipeline_bridge_s1_chipselect;
  wire             flash_ssram_pipeline_bridge_s1_debugaccess;
  wire             flash_ssram_pipeline_bridge_s1_end_xfer;
  wire             flash_ssram_pipeline_bridge_s1_endofpacket_from_sa;
  wire             flash_ssram_pipeline_bridge_s1_firsttransfer;
  wire             flash_ssram_pipeline_bridge_s1_grant_vector;
  wire             flash_ssram_pipeline_bridge_s1_in_a_read_cycle;
  wire             flash_ssram_pipeline_bridge_s1_in_a_write_cycle;
  wire             flash_ssram_pipeline_bridge_s1_master_qreq_vector;
  wire             flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction;
  wire    [ 19: 0] flash_ssram_pipeline_bridge_s1_nativeaddress;
  wire             flash_ssram_pipeline_bridge_s1_non_bursting_master_requests;
  wire             flash_ssram_pipeline_bridge_s1_read;
  wire    [255: 0] flash_ssram_pipeline_bridge_s1_readdata_from_sa;
  wire             flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa;
  reg              flash_ssram_pipeline_bridge_s1_reg_firsttransfer;
  wire             flash_ssram_pipeline_bridge_s1_reset_n;
  reg              flash_ssram_pipeline_bridge_s1_slavearbiterlockenable;
  wire             flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2;
  wire             flash_ssram_pipeline_bridge_s1_unreg_firsttransfer;
  wire             flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
  wire             flash_ssram_pipeline_bridge_s1_waits_for_read;
  wire             flash_ssram_pipeline_bridge_s1_waits_for_write;
  wire             flash_ssram_pipeline_bridge_s1_write;
  wire    [255: 0] flash_ssram_pipeline_bridge_s1_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire    [ 31: 0] pipeline_bridge_m1_byteenable_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  wire             pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_saved_grant_flash_ssram_pipeline_bridge_s1;
  wire    [255: 0] pipeline_bridge_m1_writedata_replicated;
  wire    [ 26: 0] shifted_address_to_flash_ssram_pipeline_bridge_s1_from_pipeline_bridge_m1;
  wire             wait_for_flash_ssram_pipeline_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~flash_ssram_pipeline_bridge_s1_end_xfer;
    end


  assign flash_ssram_pipeline_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1));
  //assign flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa = flash_ssram_pipeline_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa = flash_ssram_pipeline_bridge_s1_readdatavalid;

  //assign flash_ssram_pipeline_bridge_s1_readdata_from_sa = flash_ssram_pipeline_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_readdata_from_sa = flash_ssram_pipeline_bridge_s1_readdata;

  assign pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1 = ({pipeline_bridge_m1_address_to_slave[26 : 25] , 25'b0} == 27'h2000000) & pipeline_bridge_m1_chipselect;
  //assign flash_ssram_pipeline_bridge_s1_waitrequest_from_sa = flash_ssram_pipeline_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_waitrequest_from_sa = flash_ssram_pipeline_bridge_s1_waitrequest;

  //flash_ssram_pipeline_bridge_s1_arb_share_counter set values, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_arb_share_set_values = 1;

  //flash_ssram_pipeline_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_non_bursting_master_requests = pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1 |
    pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;

  //flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant = 0;

  //flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value = flash_ssram_pipeline_bridge_s1_firsttransfer ? (flash_ssram_pipeline_bridge_s1_arb_share_set_values - 1) : |flash_ssram_pipeline_bridge_s1_arb_share_counter ? (flash_ssram_pipeline_bridge_s1_arb_share_counter - 1) : 0;

  //flash_ssram_pipeline_bridge_s1_allgrants all slave grants, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_allgrants = (|flash_ssram_pipeline_bridge_s1_grant_vector) |
    (|flash_ssram_pipeline_bridge_s1_grant_vector);

  //flash_ssram_pipeline_bridge_s1_end_xfer assignment, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_end_xfer = ~(flash_ssram_pipeline_bridge_s1_waits_for_read | flash_ssram_pipeline_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 = flash_ssram_pipeline_bridge_s1_end_xfer & (~flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //flash_ssram_pipeline_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 & flash_ssram_pipeline_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 & ~flash_ssram_pipeline_bridge_s1_non_bursting_master_requests);

  //flash_ssram_pipeline_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_s1_arb_share_counter <= 0;
      else if (flash_ssram_pipeline_bridge_s1_arb_counter_enable)
          flash_ssram_pipeline_bridge_s1_arb_share_counter <= flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //flash_ssram_pipeline_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|flash_ssram_pipeline_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1) | (end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 & ~flash_ssram_pipeline_bridge_s1_non_bursting_master_requests))
          flash_ssram_pipeline_bridge_s1_slavearbiterlockenable <= |flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 flash_ssram_pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = flash_ssram_pipeline_bridge_s1_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 = |flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;

  //pipeline_bridge/m1 flash_ssram_pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //flash_ssram_pipeline_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1 = pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1 & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0) | (1 < pipeline_bridge_m1_latency_counter) | (|pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register))));
  //unique name for flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction = flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_pipeline_bridge_m1_to_flash_ssram_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pipeline_bridge_m1_to_flash_ssram_pipeline_bridge_s1_module rdv_fifo_for_pipeline_bridge_m1_to_flash_ssram_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1),
      .data_out             (pipeline_bridge_m1_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (pipeline_bridge_m1_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1),
      .full                 (),
      .read                 (flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~flash_ssram_pipeline_bridge_s1_waits_for_read)
    );

  assign pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register = ~pipeline_bridge_m1_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1;
  //local readdatavalid pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1 = flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa;

  //replicate narrow data for wide slave
  assign pipeline_bridge_m1_writedata_replicated = {pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata,
    pipeline_bridge_m1_writedata};

  //flash_ssram_pipeline_bridge_s1_writedata mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_writedata = pipeline_bridge_m1_writedata_replicated;

  //assign flash_ssram_pipeline_bridge_s1_endofpacket_from_sa = flash_ssram_pipeline_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_endofpacket_from_sa = flash_ssram_pipeline_bridge_s1_endofpacket;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1 = pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1;

  //pipeline_bridge/m1 saved-grant flash_ssram_pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_flash_ssram_pipeline_bridge_s1 = pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;

  //allow new arb cycle for flash_ssram_pipeline_bridge/s1, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign flash_ssram_pipeline_bridge_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign flash_ssram_pipeline_bridge_s1_master_qreq_vector = 1;

  //flash_ssram_pipeline_bridge_s1_reset_n assignment, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_reset_n = reset_n;

  assign flash_ssram_pipeline_bridge_s1_chipselect = pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1;
  //flash_ssram_pipeline_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_firsttransfer = flash_ssram_pipeline_bridge_s1_begins_xfer ? flash_ssram_pipeline_bridge_s1_unreg_firsttransfer : flash_ssram_pipeline_bridge_s1_reg_firsttransfer;

  //flash_ssram_pipeline_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_unreg_firsttransfer = ~(flash_ssram_pipeline_bridge_s1_slavearbiterlockenable & flash_ssram_pipeline_bridge_s1_any_continuerequest);

  //flash_ssram_pipeline_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (flash_ssram_pipeline_bridge_s1_begins_xfer)
          flash_ssram_pipeline_bridge_s1_reg_firsttransfer <= flash_ssram_pipeline_bridge_s1_unreg_firsttransfer;
    end


  //flash_ssram_pipeline_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_beginbursttransfer_internal = flash_ssram_pipeline_bridge_s1_begins_xfer;

  //flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal = flash_ssram_pipeline_bridge_s1_begins_xfer & flash_ssram_pipeline_bridge_s1_firsttransfer;

  //flash_ssram_pipeline_bridge_s1_read assignment, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_read = pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //flash_ssram_pipeline_bridge_s1_write assignment, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_write = pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_flash_ssram_pipeline_bridge_s1_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //flash_ssram_pipeline_bridge_s1_address mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_address = shifted_address_to_flash_ssram_pipeline_bridge_s1_from_pipeline_bridge_m1 >> 5;

  //slaveid flash_ssram_pipeline_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_nativeaddress = pipeline_bridge_m1_address_to_slave >> 2;

  //d1_flash_ssram_pipeline_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_flash_ssram_pipeline_bridge_s1_end_xfer <= 1;
      else 
        d1_flash_ssram_pipeline_bridge_s1_end_xfer <= flash_ssram_pipeline_bridge_s1_end_xfer;
    end


  //flash_ssram_pipeline_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_waits_for_read = flash_ssram_pipeline_bridge_s1_in_a_read_cycle & flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;

  //flash_ssram_pipeline_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_in_a_read_cycle = pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = flash_ssram_pipeline_bridge_s1_in_a_read_cycle;

  //flash_ssram_pipeline_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_waits_for_write = flash_ssram_pipeline_bridge_s1_in_a_write_cycle & flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;

  //flash_ssram_pipeline_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign flash_ssram_pipeline_bridge_s1_in_a_write_cycle = pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = flash_ssram_pipeline_bridge_s1_in_a_write_cycle;

  assign wait_for_flash_ssram_pipeline_bridge_s1_counter = 0;
  //flash_ssram_pipeline_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_byteenable = (pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1)? pipeline_bridge_m1_byteenable_flash_ssram_pipeline_bridge_s1 :
    -1;

  //byte_enable_mux for pipeline_bridge/m1 and flash_ssram_pipeline_bridge/s1, which is an e_mux
  assign pipeline_bridge_m1_byteenable_flash_ssram_pipeline_bridge_s1 = (pipeline_bridge_m1_address_to_slave[4 : 2] == 0)? pipeline_bridge_m1_byteenable :
    (pipeline_bridge_m1_address_to_slave[4 : 2] == 1)? {pipeline_bridge_m1_byteenable, {4'b0}} :
    (pipeline_bridge_m1_address_to_slave[4 : 2] == 2)? {pipeline_bridge_m1_byteenable, {8'b0}} :
    (pipeline_bridge_m1_address_to_slave[4 : 2] == 3)? {pipeline_bridge_m1_byteenable, {12'b0}} :
    (pipeline_bridge_m1_address_to_slave[4 : 2] == 4)? {pipeline_bridge_m1_byteenable, {16'b0}} :
    (pipeline_bridge_m1_address_to_slave[4 : 2] == 5)? {pipeline_bridge_m1_byteenable, {20'b0}} :
    (pipeline_bridge_m1_address_to_slave[4 : 2] == 6)? {pipeline_bridge_m1_byteenable, {24'b0}} :
    {pipeline_bridge_m1_byteenable, {28'b0}};

  //burstcount mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_burstcount = (pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1)? pipeline_bridge_m1_burstcount :
    1;

  //flash_ssram_pipeline_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_arbiterlock = pipeline_bridge_m1_arbiterlock;

  //flash_ssram_pipeline_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_arbiterlock2 = pipeline_bridge_m1_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_s1_debugaccess = (pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1)? pipeline_bridge_m1_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //flash_ssram_pipeline_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1 && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave flash_ssram_pipeline_bridge/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_ssram_pipeline_bridge_m1_arbitrator (
                                                   // inputs:
                                                    clk,
                                                    d1_tristate_bridge_avalon_slave_end_xfer,
                                                    flash_s1_wait_counter_eq_0,
                                                    flash_ssram_pipeline_bridge_m1_address,
                                                    flash_ssram_pipeline_bridge_m1_burstcount,
                                                    flash_ssram_pipeline_bridge_m1_byteenable,
                                                    flash_ssram_pipeline_bridge_m1_byteenable_flash_s1,
                                                    flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1,
                                                    flash_ssram_pipeline_bridge_m1_chipselect,
                                                    flash_ssram_pipeline_bridge_m1_granted_flash_s1,
                                                    flash_ssram_pipeline_bridge_m1_granted_ssram_s1,
                                                    flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1,
                                                    flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1,
                                                    flash_ssram_pipeline_bridge_m1_read,
                                                    flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1,
                                                    flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1,
                                                    flash_ssram_pipeline_bridge_m1_requests_flash_s1,
                                                    flash_ssram_pipeline_bridge_m1_requests_ssram_s1,
                                                    flash_ssram_pipeline_bridge_m1_write,
                                                    flash_ssram_pipeline_bridge_m1_writedata,
                                                    incoming_tristate_bridge_data,
                                                    incoming_tristate_bridge_data_with_Xs_converted_to_0,
                                                    reset_n,

                                                   // outputs:
                                                    flash_ssram_pipeline_bridge_m1_address_to_slave,
                                                    flash_ssram_pipeline_bridge_m1_dbs_address,
                                                    flash_ssram_pipeline_bridge_m1_dbs_write_16,
                                                    flash_ssram_pipeline_bridge_m1_dbs_write_32,
                                                    flash_ssram_pipeline_bridge_m1_latency_counter,
                                                    flash_ssram_pipeline_bridge_m1_readdata,
                                                    flash_ssram_pipeline_bridge_m1_readdatavalid,
                                                    flash_ssram_pipeline_bridge_m1_waitrequest
                                                 )
;

  output  [ 24: 0] flash_ssram_pipeline_bridge_m1_address_to_slave;
  output  [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_address;
  output  [ 15: 0] flash_ssram_pipeline_bridge_m1_dbs_write_16;
  output  [ 31: 0] flash_ssram_pipeline_bridge_m1_dbs_write_32;
  output  [  2: 0] flash_ssram_pipeline_bridge_m1_latency_counter;
  output  [255: 0] flash_ssram_pipeline_bridge_m1_readdata;
  output           flash_ssram_pipeline_bridge_m1_readdatavalid;
  output           flash_ssram_pipeline_bridge_m1_waitrequest;
  input            clk;
  input            d1_tristate_bridge_avalon_slave_end_xfer;
  input            flash_s1_wait_counter_eq_0;
  input   [ 24: 0] flash_ssram_pipeline_bridge_m1_address;
  input            flash_ssram_pipeline_bridge_m1_burstcount;
  input   [ 31: 0] flash_ssram_pipeline_bridge_m1_byteenable;
  input   [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1;
  input   [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1;
  input            flash_ssram_pipeline_bridge_m1_chipselect;
  input            flash_ssram_pipeline_bridge_m1_granted_flash_s1;
  input            flash_ssram_pipeline_bridge_m1_granted_ssram_s1;
  input            flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1;
  input            flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1;
  input            flash_ssram_pipeline_bridge_m1_read;
  input            flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1;
  input            flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1;
  input            flash_ssram_pipeline_bridge_m1_requests_flash_s1;
  input            flash_ssram_pipeline_bridge_m1_requests_ssram_s1;
  input            flash_ssram_pipeline_bridge_m1_write;
  input   [255: 0] flash_ssram_pipeline_bridge_m1_writedata;
  input   [ 31: 0] incoming_tristate_bridge_data;
  input   [ 15: 0] incoming_tristate_bridge_data_with_Xs_converted_to_0;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  reg     [ 15: 0] dbs_latent_16_reg_segment_1;
  reg     [ 15: 0] dbs_latent_16_reg_segment_10;
  reg     [ 15: 0] dbs_latent_16_reg_segment_11;
  reg     [ 15: 0] dbs_latent_16_reg_segment_12;
  reg     [ 15: 0] dbs_latent_16_reg_segment_13;
  reg     [ 15: 0] dbs_latent_16_reg_segment_14;
  reg     [ 15: 0] dbs_latent_16_reg_segment_2;
  reg     [ 15: 0] dbs_latent_16_reg_segment_3;
  reg     [ 15: 0] dbs_latent_16_reg_segment_4;
  reg     [ 15: 0] dbs_latent_16_reg_segment_5;
  reg     [ 15: 0] dbs_latent_16_reg_segment_6;
  reg     [ 15: 0] dbs_latent_16_reg_segment_7;
  reg     [ 15: 0] dbs_latent_16_reg_segment_8;
  reg     [ 15: 0] dbs_latent_16_reg_segment_9;
  reg     [ 31: 0] dbs_latent_32_reg_segment_0;
  reg     [ 31: 0] dbs_latent_32_reg_segment_1;
  reg     [ 31: 0] dbs_latent_32_reg_segment_2;
  reg     [ 31: 0] dbs_latent_32_reg_segment_3;
  reg     [ 31: 0] dbs_latent_32_reg_segment_4;
  reg     [ 31: 0] dbs_latent_32_reg_segment_5;
  reg     [ 31: 0] dbs_latent_32_reg_segment_6;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  reg     [ 24: 0] flash_ssram_pipeline_bridge_m1_address_last_time;
  wire    [ 24: 0] flash_ssram_pipeline_bridge_m1_address_to_slave;
  reg              flash_ssram_pipeline_bridge_m1_burstcount_last_time;
  reg     [ 31: 0] flash_ssram_pipeline_bridge_m1_byteenable_last_time;
  reg              flash_ssram_pipeline_bridge_m1_chipselect_last_time;
  reg     [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_address;
  wire    [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_increment;
  reg     [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_rdv_counter;
  wire    [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_rdv_counter_inc;
  wire    [ 15: 0] flash_ssram_pipeline_bridge_m1_dbs_write_16;
  wire    [ 31: 0] flash_ssram_pipeline_bridge_m1_dbs_write_32;
  wire             flash_ssram_pipeline_bridge_m1_is_granted_some_slave;
  reg     [  2: 0] flash_ssram_pipeline_bridge_m1_latency_counter;
  wire    [  4: 0] flash_ssram_pipeline_bridge_m1_next_dbs_rdv_counter;
  reg              flash_ssram_pipeline_bridge_m1_read_but_no_slave_selected;
  reg              flash_ssram_pipeline_bridge_m1_read_last_time;
  wire    [255: 0] flash_ssram_pipeline_bridge_m1_readdata;
  wire             flash_ssram_pipeline_bridge_m1_readdatavalid;
  wire             flash_ssram_pipeline_bridge_m1_run;
  wire             flash_ssram_pipeline_bridge_m1_waitrequest;
  reg              flash_ssram_pipeline_bridge_m1_write_last_time;
  reg     [255: 0] flash_ssram_pipeline_bridge_m1_writedata_last_time;
  wire    [  2: 0] latency_load_value;
  wire    [  4: 0] next_dbs_address;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_1;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_10;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_11;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_12;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_13;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_14;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_2;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_3;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_4;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_5;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_6;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_7;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_8;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_9;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_0;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_1;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_2;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_3;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_4;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_5;
  wire    [ 31: 0] p1_dbs_latent_32_reg_segment_6;
  wire    [  2: 0] p1_flash_ssram_pipeline_bridge_m1_latency_counter;
  wire             pre_dbs_count_enable;
  wire             pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & ((flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 | (((flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) & !flash_ssram_pipeline_bridge_m1_byteenable_flash_s1 & flash_ssram_pipeline_bridge_m1_dbs_address[4] & flash_ssram_pipeline_bridge_m1_dbs_address[3] & flash_ssram_pipeline_bridge_m1_dbs_address[2] & flash_ssram_pipeline_bridge_m1_dbs_address[1])) | ~flash_ssram_pipeline_bridge_m1_requests_flash_s1)) & ((flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1 | (((flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) & !flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1 & flash_ssram_pipeline_bridge_m1_dbs_address[4] & flash_ssram_pipeline_bridge_m1_dbs_address[3] & flash_ssram_pipeline_bridge_m1_dbs_address[2])) | ~flash_ssram_pipeline_bridge_m1_requests_ssram_s1)) & ((~flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 | ~(flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) | (1 & ((flash_s1_wait_counter_eq_0 & ~d1_tristate_bridge_avalon_slave_end_xfer)) & (flash_ssram_pipeline_bridge_m1_dbs_address[4] & flash_ssram_pipeline_bridge_m1_dbs_address[3] & flash_ssram_pipeline_bridge_m1_dbs_address[2] & flash_ssram_pipeline_bridge_m1_dbs_address[1]) & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect)))) & ((~flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 | ~(flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) | (1 & ((flash_s1_wait_counter_eq_0 & ~d1_tristate_bridge_avalon_slave_end_xfer)) & (flash_ssram_pipeline_bridge_m1_dbs_address[4] & flash_ssram_pipeline_bridge_m1_dbs_address[3] & flash_ssram_pipeline_bridge_m1_dbs_address[2] & flash_ssram_pipeline_bridge_m1_dbs_address[1]) & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect)))) & ((~flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1 | ~(flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) | (1 & (flash_ssram_pipeline_bridge_m1_dbs_address[4] & flash_ssram_pipeline_bridge_m1_dbs_address[3] & flash_ssram_pipeline_bridge_m1_dbs_address[2]) & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect)))) & ((~flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1 | ~(flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) | (1 & (flash_ssram_pipeline_bridge_m1_dbs_address[4] & flash_ssram_pipeline_bridge_m1_dbs_address[3] & flash_ssram_pipeline_bridge_m1_dbs_address[2]) & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect))));

  //cascaded wait assignment, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign flash_ssram_pipeline_bridge_m1_address_to_slave = flash_ssram_pipeline_bridge_m1_address[24 : 0];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & flash_ssram_pipeline_bridge_m1_requests_flash_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) & !flash_ssram_pipeline_bridge_m1_byteenable_flash_s1)) |
    (((~0) & flash_ssram_pipeline_bridge_m1_requests_ssram_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) & !flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1)) |
    ((flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & 1 & 1 & ({flash_s1_wait_counter_eq_0 & ~d1_tristate_bridge_avalon_slave_end_xfer}))) |
    ((flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) & 1 & 1 & ({flash_s1_wait_counter_eq_0 & ~d1_tristate_bridge_avalon_slave_end_xfer}))) |
    ((flash_ssram_pipeline_bridge_m1_granted_ssram_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & 1 & 1)) |
    ((flash_ssram_pipeline_bridge_m1_granted_ssram_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect) & 1 & 1));

  //flash_ssram_pipeline_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_read_but_no_slave_selected <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_read_but_no_slave_selected <= (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & flash_ssram_pipeline_bridge_m1_run & ~flash_ssram_pipeline_bridge_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_is_granted_some_slave = flash_ssram_pipeline_bridge_m1_granted_flash_s1 |
    flash_ssram_pipeline_bridge_m1_granted_ssram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid = (flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1 & dbs_rdv_counter_overflow) |
    (flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1 & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_readdatavalid = flash_ssram_pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid |
    flash_ssram_pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid;

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //input to latent dbs-16 stored 1, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_1 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_1 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 1))
          dbs_latent_16_reg_segment_1 <= p1_dbs_latent_16_reg_segment_1;
    end


  //input to latent dbs-16 stored 2, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_2 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_2 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 2))
          dbs_latent_16_reg_segment_2 <= p1_dbs_latent_16_reg_segment_2;
    end


  //input to latent dbs-16 stored 3, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_3 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_3 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 3))
          dbs_latent_16_reg_segment_3 <= p1_dbs_latent_16_reg_segment_3;
    end


  //input to latent dbs-16 stored 4, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_4 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_4 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 4))
          dbs_latent_16_reg_segment_4 <= p1_dbs_latent_16_reg_segment_4;
    end


  //input to latent dbs-16 stored 5, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_5 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_5 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 5))
          dbs_latent_16_reg_segment_5 <= p1_dbs_latent_16_reg_segment_5;
    end


  //input to latent dbs-16 stored 6, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_6 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_6 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 6))
          dbs_latent_16_reg_segment_6 <= p1_dbs_latent_16_reg_segment_6;
    end


  //input to latent dbs-16 stored 7, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_7 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_7 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 7))
          dbs_latent_16_reg_segment_7 <= p1_dbs_latent_16_reg_segment_7;
    end


  //input to latent dbs-16 stored 8, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_8 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_8 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 8))
          dbs_latent_16_reg_segment_8 <= p1_dbs_latent_16_reg_segment_8;
    end


  //input to latent dbs-16 stored 9, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_9 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_9 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 9))
          dbs_latent_16_reg_segment_9 <= p1_dbs_latent_16_reg_segment_9;
    end


  //input to latent dbs-16 stored 10, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_10 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_10 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 10))
          dbs_latent_16_reg_segment_10 <= p1_dbs_latent_16_reg_segment_10;
    end


  //input to latent dbs-16 stored 11, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_11 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_11 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 11))
          dbs_latent_16_reg_segment_11 <= p1_dbs_latent_16_reg_segment_11;
    end


  //input to latent dbs-16 stored 12, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_12 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_12 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 12))
          dbs_latent_16_reg_segment_12 <= p1_dbs_latent_16_reg_segment_12;
    end


  //input to latent dbs-16 stored 13, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_13 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_13 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 13))
          dbs_latent_16_reg_segment_13 <= p1_dbs_latent_16_reg_segment_13;
    end


  //input to latent dbs-16 stored 14, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_14 = incoming_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_14 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 1]) == 14))
          dbs_latent_16_reg_segment_14 <= p1_dbs_latent_16_reg_segment_14;
    end


  //flash_ssram_pipeline_bridge/m1 readdata mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_readdata = ({256 {~flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1}} | {incoming_tristate_bridge_data_with_Xs_converted_to_0[15 : 0],
    dbs_latent_16_reg_segment_14,
    dbs_latent_16_reg_segment_13,
    dbs_latent_16_reg_segment_12,
    dbs_latent_16_reg_segment_11,
    dbs_latent_16_reg_segment_10,
    dbs_latent_16_reg_segment_9,
    dbs_latent_16_reg_segment_8,
    dbs_latent_16_reg_segment_7,
    dbs_latent_16_reg_segment_6,
    dbs_latent_16_reg_segment_5,
    dbs_latent_16_reg_segment_4,
    dbs_latent_16_reg_segment_3,
    dbs_latent_16_reg_segment_2,
    dbs_latent_16_reg_segment_1,
    dbs_latent_16_reg_segment_0}) &
    ({256 {~flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1}} | {incoming_tristate_bridge_data[31 : 0],
    dbs_latent_32_reg_segment_6,
    dbs_latent_32_reg_segment_5,
    dbs_latent_32_reg_segment_4,
    dbs_latent_32_reg_segment_3,
    dbs_latent_32_reg_segment_2,
    dbs_latent_32_reg_segment_1,
    dbs_latent_32_reg_segment_0});

  //mux write dbs 4, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_dbs_write_16 = ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 0))? flash_ssram_pipeline_bridge_m1_writedata[15 : 0] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 1))? flash_ssram_pipeline_bridge_m1_writedata[31 : 16] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 2))? flash_ssram_pipeline_bridge_m1_writedata[47 : 32] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 3))? flash_ssram_pipeline_bridge_m1_writedata[63 : 48] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 4))? flash_ssram_pipeline_bridge_m1_writedata[79 : 64] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 5))? flash_ssram_pipeline_bridge_m1_writedata[95 : 80] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 6))? flash_ssram_pipeline_bridge_m1_writedata[111 : 96] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 7))? flash_ssram_pipeline_bridge_m1_writedata[127 : 112] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 8))? flash_ssram_pipeline_bridge_m1_writedata[143 : 128] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 9))? flash_ssram_pipeline_bridge_m1_writedata[159 : 144] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 10))? flash_ssram_pipeline_bridge_m1_writedata[175 : 160] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 11))? flash_ssram_pipeline_bridge_m1_writedata[191 : 176] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 12))? flash_ssram_pipeline_bridge_m1_writedata[207 : 192] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 13))? flash_ssram_pipeline_bridge_m1_writedata[223 : 208] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 14))? flash_ssram_pipeline_bridge_m1_writedata[239 : 224] :
    flash_ssram_pipeline_bridge_m1_writedata[255 : 240];

  //actual waitrequest port, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_waitrequest = ~flash_ssram_pipeline_bridge_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_latency_counter <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_latency_counter <= p1_flash_ssram_pipeline_bridge_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_flash_ssram_pipeline_bridge_m1_latency_counter = ((flash_ssram_pipeline_bridge_m1_run & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect)))? latency_load_value :
    (flash_ssram_pipeline_bridge_m1_latency_counter)? flash_ssram_pipeline_bridge_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({3 {flash_ssram_pipeline_bridge_m1_requests_flash_s1}} & 2) |
    ({3 {flash_ssram_pipeline_bridge_m1_requests_ssram_s1}} & 4);

  //input to latent dbs-32 stored 0, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_0 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 0))
          dbs_latent_32_reg_segment_0 <= p1_dbs_latent_32_reg_segment_0;
    end


  //input to latent dbs-32 stored 1, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_1 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_1 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 1))
          dbs_latent_32_reg_segment_1 <= p1_dbs_latent_32_reg_segment_1;
    end


  //input to latent dbs-32 stored 2, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_2 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_2 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 2))
          dbs_latent_32_reg_segment_2 <= p1_dbs_latent_32_reg_segment_2;
    end


  //input to latent dbs-32 stored 3, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_3 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_3 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 3))
          dbs_latent_32_reg_segment_3 <= p1_dbs_latent_32_reg_segment_3;
    end


  //input to latent dbs-32 stored 4, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_4 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_4 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 4))
          dbs_latent_32_reg_segment_4 <= p1_dbs_latent_32_reg_segment_4;
    end


  //input to latent dbs-32 stored 5, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_5 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_5 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 5))
          dbs_latent_32_reg_segment_5 <= p1_dbs_latent_32_reg_segment_5;
    end


  //input to latent dbs-32 stored 6, which is an e_mux
  assign p1_dbs_latent_32_reg_segment_6 = incoming_tristate_bridge_data;

  //dbs register for latent dbs-32 segment 6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_32_reg_segment_6 <= 0;
      else if (dbs_rdv_count_enable & ((flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4 : 2]) == 6))
          dbs_latent_32_reg_segment_6 <= p1_dbs_latent_32_reg_segment_6;
    end


  //mux write dbs 3, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_dbs_write_32 = ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 0))? flash_ssram_pipeline_bridge_m1_writedata[31 : 0] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 1))? flash_ssram_pipeline_bridge_m1_writedata[63 : 32] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 2))? flash_ssram_pipeline_bridge_m1_writedata[95 : 64] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 3))? flash_ssram_pipeline_bridge_m1_writedata[127 : 96] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 4))? flash_ssram_pipeline_bridge_m1_writedata[159 : 128] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 5))? flash_ssram_pipeline_bridge_m1_writedata[191 : 160] :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 6))? flash_ssram_pipeline_bridge_m1_writedata[223 : 192] :
    flash_ssram_pipeline_bridge_m1_writedata[255 : 224];

  //dbs count increment, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_dbs_increment = (flash_ssram_pipeline_bridge_m1_requests_flash_s1)? 2 :
    (flash_ssram_pipeline_bridge_m1_requests_ssram_s1)? 4 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = flash_ssram_pipeline_bridge_m1_dbs_address[4] & !(next_dbs_address[4]);

  //next master address, which is an e_assign
  assign next_dbs_address = flash_ssram_pipeline_bridge_m1_dbs_address + flash_ssram_pipeline_bridge_m1_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_dbs_address <= 0;
      else if (dbs_count_enable)
          flash_ssram_pipeline_bridge_m1_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_next_dbs_rdv_counter = flash_ssram_pipeline_bridge_m1_dbs_rdv_counter + flash_ssram_pipeline_bridge_m1_dbs_rdv_counter_inc;

  //flash_ssram_pipeline_bridge_m1_rdv_inc_mux, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_dbs_rdv_counter_inc = (flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1)? 2 :
    4;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1 |
    flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          flash_ssram_pipeline_bridge_m1_dbs_rdv_counter <= flash_ssram_pipeline_bridge_m1_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = flash_ssram_pipeline_bridge_m1_dbs_rdv_counter[4] & ~flash_ssram_pipeline_bridge_m1_next_dbs_rdv_counter[4];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //flash_ssram_pipeline_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_address_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_address_last_time <= flash_ssram_pipeline_bridge_m1_address;
    end


  //flash_ssram_pipeline_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= flash_ssram_pipeline_bridge_m1_waitrequest & flash_ssram_pipeline_bridge_m1_chipselect;
    end


  //flash_ssram_pipeline_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_address != flash_ssram_pipeline_bridge_m1_address_last_time))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //flash_ssram_pipeline_bridge_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_chipselect_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_chipselect_last_time <= flash_ssram_pipeline_bridge_m1_chipselect;
    end


  //flash_ssram_pipeline_bridge_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_chipselect != flash_ssram_pipeline_bridge_m1_chipselect_last_time))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //flash_ssram_pipeline_bridge_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_burstcount_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_burstcount_last_time <= flash_ssram_pipeline_bridge_m1_burstcount;
    end


  //flash_ssram_pipeline_bridge_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_burstcount != flash_ssram_pipeline_bridge_m1_burstcount_last_time))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //flash_ssram_pipeline_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_byteenable_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_byteenable_last_time <= flash_ssram_pipeline_bridge_m1_byteenable;
    end


  //flash_ssram_pipeline_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_byteenable != flash_ssram_pipeline_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //flash_ssram_pipeline_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_read_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_read_last_time <= flash_ssram_pipeline_bridge_m1_read;
    end


  //flash_ssram_pipeline_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_read != flash_ssram_pipeline_bridge_m1_read_last_time))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //flash_ssram_pipeline_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_write_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_write_last_time <= flash_ssram_pipeline_bridge_m1_write;
    end


  //flash_ssram_pipeline_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_write != flash_ssram_pipeline_bridge_m1_write_last_time))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //flash_ssram_pipeline_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_writedata_last_time <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_writedata_last_time <= flash_ssram_pipeline_bridge_m1_writedata;
    end


  //flash_ssram_pipeline_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (flash_ssram_pipeline_bridge_m1_writedata != flash_ssram_pipeline_bridge_m1_writedata_last_time) & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect))
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_ssram_pipeline_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_ddr_sdram_clock_crossing_bridge_m1_to_frame_buffer_s1_module (
                                                                                   // inputs:
                                                                                    clear_fifo,
                                                                                    clk,
                                                                                    data_in,
                                                                                    read,
                                                                                    reset_n,
                                                                                    sync_reset,
                                                                                    write,

                                                                                   // outputs:
                                                                                    data_out,
                                                                                    empty,
                                                                                    fifo_contains_ones_n,
                                                                                    full
                                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module frame_buffer_s1_arbitrator (
                                    // inputs:
                                     clk,
                                     ddr_sdram_clock_crossing_bridge_m1_address_to_slave,
                                     ddr_sdram_clock_crossing_bridge_m1_byteenable,
                                     ddr_sdram_clock_crossing_bridge_m1_latency_counter,
                                     ddr_sdram_clock_crossing_bridge_m1_read,
                                     ddr_sdram_clock_crossing_bridge_m1_write,
                                     ddr_sdram_clock_crossing_bridge_m1_writedata,
                                     frame_buffer_s1_readdata,
                                     frame_buffer_s1_readdatavalid,
                                     frame_buffer_s1_resetrequest_n,
                                     frame_buffer_s1_waitrequest_n,
                                     reset_n,

                                    // outputs:
                                     d1_frame_buffer_s1_end_xfer,
                                     ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1,
                                     ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1,
                                     ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1,
                                     ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register,
                                     ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1,
                                     frame_buffer_s1_address,
                                     frame_buffer_s1_beginbursttransfer,
                                     frame_buffer_s1_burstcount,
                                     frame_buffer_s1_byteenable,
                                     frame_buffer_s1_read,
                                     frame_buffer_s1_readdata_from_sa,
                                     frame_buffer_s1_resetrequest_n_from_sa,
                                     frame_buffer_s1_waitrequest_n_from_sa,
                                     frame_buffer_s1_write,
                                     frame_buffer_s1_writedata
                                  )
;

  output           d1_frame_buffer_s1_end_xfer;
  output           ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1;
  output           ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1;
  output           ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1;
  output           ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register;
  output           ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1;
  output  [ 22: 0] frame_buffer_s1_address;
  output           frame_buffer_s1_beginbursttransfer;
  output  [  1: 0] frame_buffer_s1_burstcount;
  output  [  3: 0] frame_buffer_s1_byteenable;
  output           frame_buffer_s1_read;
  output  [ 31: 0] frame_buffer_s1_readdata_from_sa;
  output           frame_buffer_s1_resetrequest_n_from_sa;
  output           frame_buffer_s1_waitrequest_n_from_sa;
  output           frame_buffer_s1_write;
  output  [ 31: 0] frame_buffer_s1_writedata;
  input            clk;
  input   [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address_to_slave;
  input   [  3: 0] ddr_sdram_clock_crossing_bridge_m1_byteenable;
  input            ddr_sdram_clock_crossing_bridge_m1_latency_counter;
  input            ddr_sdram_clock_crossing_bridge_m1_read;
  input            ddr_sdram_clock_crossing_bridge_m1_write;
  input   [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] frame_buffer_s1_readdata;
  input            frame_buffer_s1_readdatavalid;
  input            frame_buffer_s1_resetrequest_n;
  input            frame_buffer_s1_waitrequest_n;
  input            reset_n;

  reg              d1_frame_buffer_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire             ddr_sdram_clock_crossing_bridge_m1_arbiterlock;
  wire             ddr_sdram_clock_crossing_bridge_m1_arbiterlock2;
  wire             ddr_sdram_clock_crossing_bridge_m1_continuerequest;
  wire             ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_rdv_fifo_empty_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_rdv_fifo_output_from_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register;
  wire             ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_saved_grant_frame_buffer_s1;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_frame_buffer_s1;
  wire    [ 22: 0] frame_buffer_s1_address;
  wire             frame_buffer_s1_allgrants;
  wire             frame_buffer_s1_allow_new_arb_cycle;
  wire             frame_buffer_s1_any_bursting_master_saved_grant;
  wire             frame_buffer_s1_any_continuerequest;
  wire             frame_buffer_s1_arb_counter_enable;
  reg              frame_buffer_s1_arb_share_counter;
  wire             frame_buffer_s1_arb_share_counter_next_value;
  wire             frame_buffer_s1_arb_share_set_values;
  reg              frame_buffer_s1_bbt_burstcounter;
  wire             frame_buffer_s1_beginbursttransfer;
  wire             frame_buffer_s1_beginbursttransfer_internal;
  wire             frame_buffer_s1_begins_xfer;
  wire    [  1: 0] frame_buffer_s1_burstcount;
  wire    [  3: 0] frame_buffer_s1_byteenable;
  wire             frame_buffer_s1_end_xfer;
  wire             frame_buffer_s1_firsttransfer;
  wire             frame_buffer_s1_grant_vector;
  wire             frame_buffer_s1_in_a_read_cycle;
  wire             frame_buffer_s1_in_a_write_cycle;
  wire             frame_buffer_s1_master_qreq_vector;
  wire             frame_buffer_s1_move_on_to_next_transaction;
  wire             frame_buffer_s1_next_bbt_burstcount;
  wire             frame_buffer_s1_non_bursting_master_requests;
  wire             frame_buffer_s1_read;
  wire    [ 31: 0] frame_buffer_s1_readdata_from_sa;
  wire             frame_buffer_s1_readdatavalid_from_sa;
  reg              frame_buffer_s1_reg_firsttransfer;
  wire             frame_buffer_s1_resetrequest_n_from_sa;
  reg              frame_buffer_s1_slavearbiterlockenable;
  wire             frame_buffer_s1_slavearbiterlockenable2;
  wire             frame_buffer_s1_unreg_firsttransfer;
  wire             frame_buffer_s1_waitrequest_n_from_sa;
  wire             frame_buffer_s1_waits_for_read;
  wire             frame_buffer_s1_waits_for_write;
  wire             frame_buffer_s1_write;
  wire    [ 31: 0] frame_buffer_s1_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 24: 0] shifted_address_to_frame_buffer_s1_from_ddr_sdram_clock_crossing_bridge_m1;
  wire             wait_for_frame_buffer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~frame_buffer_s1_end_xfer;
    end


  assign frame_buffer_s1_begins_xfer = ~d1_reasons_to_wait & ((ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1));
  //assign frame_buffer_s1_readdata_from_sa = frame_buffer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_s1_readdata_from_sa = frame_buffer_s1_readdata;

  assign ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1 = (1) & (ddr_sdram_clock_crossing_bridge_m1_read | ddr_sdram_clock_crossing_bridge_m1_write);
  //assign frame_buffer_s1_waitrequest_n_from_sa = frame_buffer_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_s1_waitrequest_n_from_sa = frame_buffer_s1_waitrequest_n;

  //assign frame_buffer_s1_readdatavalid_from_sa = frame_buffer_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_s1_readdatavalid_from_sa = frame_buffer_s1_readdatavalid;

  //frame_buffer_s1_arb_share_counter set values, which is an e_mux
  assign frame_buffer_s1_arb_share_set_values = 1;

  //frame_buffer_s1_non_bursting_master_requests mux, which is an e_mux
  assign frame_buffer_s1_non_bursting_master_requests = ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1;

  //frame_buffer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign frame_buffer_s1_any_bursting_master_saved_grant = 0;

  //frame_buffer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign frame_buffer_s1_arb_share_counter_next_value = frame_buffer_s1_firsttransfer ? (frame_buffer_s1_arb_share_set_values - 1) : |frame_buffer_s1_arb_share_counter ? (frame_buffer_s1_arb_share_counter - 1) : 0;

  //frame_buffer_s1_allgrants all slave grants, which is an e_mux
  assign frame_buffer_s1_allgrants = |frame_buffer_s1_grant_vector;

  //frame_buffer_s1_end_xfer assignment, which is an e_assign
  assign frame_buffer_s1_end_xfer = ~(frame_buffer_s1_waits_for_read | frame_buffer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_frame_buffer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_frame_buffer_s1 = frame_buffer_s1_end_xfer & (~frame_buffer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //frame_buffer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign frame_buffer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_frame_buffer_s1 & frame_buffer_s1_allgrants) | (end_xfer_arb_share_counter_term_frame_buffer_s1 & ~frame_buffer_s1_non_bursting_master_requests);

  //frame_buffer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_s1_arb_share_counter <= 0;
      else if (frame_buffer_s1_arb_counter_enable)
          frame_buffer_s1_arb_share_counter <= frame_buffer_s1_arb_share_counter_next_value;
    end


  //frame_buffer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_s1_slavearbiterlockenable <= 0;
      else if ((|frame_buffer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_frame_buffer_s1) | (end_xfer_arb_share_counter_term_frame_buffer_s1 & ~frame_buffer_s1_non_bursting_master_requests))
          frame_buffer_s1_slavearbiterlockenable <= |frame_buffer_s1_arb_share_counter_next_value;
    end


  //ddr_sdram_clock_crossing_bridge/m1 frame_buffer/s1 arbiterlock, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_arbiterlock = frame_buffer_s1_slavearbiterlockenable & ddr_sdram_clock_crossing_bridge_m1_continuerequest;

  //frame_buffer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign frame_buffer_s1_slavearbiterlockenable2 = |frame_buffer_s1_arb_share_counter_next_value;

  //ddr_sdram_clock_crossing_bridge/m1 frame_buffer/s1 arbiterlock2, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_arbiterlock2 = frame_buffer_s1_slavearbiterlockenable2 & ddr_sdram_clock_crossing_bridge_m1_continuerequest;

  //frame_buffer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign frame_buffer_s1_any_continuerequest = 1;

  //ddr_sdram_clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_continuerequest = 1;

  assign ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1 = ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1 & ~((ddr_sdram_clock_crossing_bridge_m1_read & ((ddr_sdram_clock_crossing_bridge_m1_latency_counter != 0) | (1 < ddr_sdram_clock_crossing_bridge_m1_latency_counter))));
  //unique name for frame_buffer_s1_move_on_to_next_transaction, which is an e_assign
  assign frame_buffer_s1_move_on_to_next_transaction = frame_buffer_s1_readdatavalid_from_sa;

  //rdv_fifo_for_ddr_sdram_clock_crossing_bridge_m1_to_frame_buffer_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_ddr_sdram_clock_crossing_bridge_m1_to_frame_buffer_s1_module rdv_fifo_for_ddr_sdram_clock_crossing_bridge_m1_to_frame_buffer_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1),
      .data_out             (ddr_sdram_clock_crossing_bridge_m1_rdv_fifo_output_from_frame_buffer_s1),
      .empty                (),
      .fifo_contains_ones_n (ddr_sdram_clock_crossing_bridge_m1_rdv_fifo_empty_frame_buffer_s1),
      .full                 (),
      .read                 (frame_buffer_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~frame_buffer_s1_waits_for_read)
    );

  assign ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register = ~ddr_sdram_clock_crossing_bridge_m1_rdv_fifo_empty_frame_buffer_s1;
  //local readdatavalid ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1, which is an e_mux
  assign ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1 = frame_buffer_s1_readdatavalid_from_sa;

  //frame_buffer_s1_writedata mux, which is an e_mux
  assign frame_buffer_s1_writedata = ddr_sdram_clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1 = ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1;

  //ddr_sdram_clock_crossing_bridge/m1 saved-grant frame_buffer/s1, which is an e_assign
  assign ddr_sdram_clock_crossing_bridge_m1_saved_grant_frame_buffer_s1 = ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1;

  //allow new arb cycle for frame_buffer/s1, which is an e_assign
  assign frame_buffer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign frame_buffer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign frame_buffer_s1_master_qreq_vector = 1;

  //assign frame_buffer_s1_resetrequest_n_from_sa = frame_buffer_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_s1_resetrequest_n_from_sa = frame_buffer_s1_resetrequest_n;

  //frame_buffer_s1_firsttransfer first transaction, which is an e_assign
  assign frame_buffer_s1_firsttransfer = frame_buffer_s1_begins_xfer ? frame_buffer_s1_unreg_firsttransfer : frame_buffer_s1_reg_firsttransfer;

  //frame_buffer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign frame_buffer_s1_unreg_firsttransfer = ~(frame_buffer_s1_slavearbiterlockenable & frame_buffer_s1_any_continuerequest);

  //frame_buffer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_s1_reg_firsttransfer <= 1'b1;
      else if (frame_buffer_s1_begins_xfer)
          frame_buffer_s1_reg_firsttransfer <= frame_buffer_s1_unreg_firsttransfer;
    end


  //frame_buffer_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign frame_buffer_s1_next_bbt_burstcount = ((((frame_buffer_s1_write) && (frame_buffer_s1_bbt_burstcounter == 0))))? (frame_buffer_s1_burstcount - 1) :
    ((((frame_buffer_s1_read) && (frame_buffer_s1_bbt_burstcounter == 0))))? 0 :
    (frame_buffer_s1_bbt_burstcounter - 1);

  //frame_buffer_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_s1_bbt_burstcounter <= 0;
      else if (frame_buffer_s1_begins_xfer)
          frame_buffer_s1_bbt_burstcounter <= frame_buffer_s1_next_bbt_burstcount;
    end


  //frame_buffer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign frame_buffer_s1_beginbursttransfer_internal = frame_buffer_s1_begins_xfer & (frame_buffer_s1_bbt_burstcounter == 0);

  //frame_buffer/s1 begin burst transfer to slave, which is an e_assign
  assign frame_buffer_s1_beginbursttransfer = frame_buffer_s1_beginbursttransfer_internal;

  //frame_buffer_s1_read assignment, which is an e_mux
  assign frame_buffer_s1_read = ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1 & ddr_sdram_clock_crossing_bridge_m1_read;

  //frame_buffer_s1_write assignment, which is an e_mux
  assign frame_buffer_s1_write = ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1 & ddr_sdram_clock_crossing_bridge_m1_write;

  assign shifted_address_to_frame_buffer_s1_from_ddr_sdram_clock_crossing_bridge_m1 = ddr_sdram_clock_crossing_bridge_m1_address_to_slave;
  //frame_buffer_s1_address mux, which is an e_mux
  assign frame_buffer_s1_address = shifted_address_to_frame_buffer_s1_from_ddr_sdram_clock_crossing_bridge_m1 >> 2;

  //d1_frame_buffer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_frame_buffer_s1_end_xfer <= 1;
      else 
        d1_frame_buffer_s1_end_xfer <= frame_buffer_s1_end_xfer;
    end


  //frame_buffer_s1_waits_for_read in a cycle, which is an e_mux
  assign frame_buffer_s1_waits_for_read = frame_buffer_s1_in_a_read_cycle & ~frame_buffer_s1_waitrequest_n_from_sa;

  //frame_buffer_s1_in_a_read_cycle assignment, which is an e_assign
  assign frame_buffer_s1_in_a_read_cycle = ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1 & ddr_sdram_clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = frame_buffer_s1_in_a_read_cycle;

  //frame_buffer_s1_waits_for_write in a cycle, which is an e_mux
  assign frame_buffer_s1_waits_for_write = frame_buffer_s1_in_a_write_cycle & ~frame_buffer_s1_waitrequest_n_from_sa;

  //frame_buffer_s1_in_a_write_cycle assignment, which is an e_assign
  assign frame_buffer_s1_in_a_write_cycle = ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1 & ddr_sdram_clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = frame_buffer_s1_in_a_write_cycle;

  assign wait_for_frame_buffer_s1_counter = 0;
  //frame_buffer_s1_byteenable byte enable port mux, which is an e_mux
  assign frame_buffer_s1_byteenable = (ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1)? ddr_sdram_clock_crossing_bridge_m1_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign frame_buffer_s1_burstcount = 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //frame_buffer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_reset_ext_clk_one_domain_synch_module (
                                                      // inputs:
                                                       clk,
                                                       data_in,
                                                       reset_n,

                                                      // outputs:
                                                       data_out
                                                    )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_lcd_sgdma_m_read_to_frame_buffer_pipeline_bridge_s1_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  wire             full_51;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_50;
  assign empty = !full_0;
  assign full_51 = 0;
  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    0;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_pipeline_bridge_m1_to_frame_buffer_pipeline_bridge_s1_module (
                                                                                   // inputs:
                                                                                    clear_fifo,
                                                                                    clk,
                                                                                    data_in,
                                                                                    read,
                                                                                    reset_n,
                                                                                    sync_reset,
                                                                                    write,

                                                                                   // outputs:
                                                                                    data_out,
                                                                                    empty,
                                                                                    fifo_contains_ones_n,
                                                                                    full
                                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  wire             full_51;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_50;
  assign empty = !full_0;
  assign full_51 = 0;
  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    0;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module frame_buffer_pipeline_bridge_s1_arbitrator (
                                                    // inputs:
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave,
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable,
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write,
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata,
                                                     clk,
                                                     frame_buffer_pipeline_bridge_s1_endofpacket,
                                                     frame_buffer_pipeline_bridge_s1_readdata,
                                                     frame_buffer_pipeline_bridge_s1_readdatavalid,
                                                     frame_buffer_pipeline_bridge_s1_waitrequest,
                                                     lcd_sgdma_m_read_address_to_slave,
                                                     lcd_sgdma_m_read_latency_counter,
                                                     lcd_sgdma_m_read_read,
                                                     pipeline_bridge_m1_address_to_slave,
                                                     pipeline_bridge_m1_burstcount,
                                                     pipeline_bridge_m1_byteenable,
                                                     pipeline_bridge_m1_chipselect,
                                                     pipeline_bridge_m1_debugaccess,
                                                     pipeline_bridge_m1_latency_counter,
                                                     pipeline_bridge_m1_read,
                                                     pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                                     pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                                     pipeline_bridge_m1_write,
                                                     pipeline_bridge_m1_writedata,
                                                     reset_n,

                                                    // outputs:
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1,
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1,
                                                     accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1,
                                                     d1_frame_buffer_pipeline_bridge_s1_end_xfer,
                                                     frame_buffer_pipeline_bridge_s1_address,
                                                     frame_buffer_pipeline_bridge_s1_arbiterlock,
                                                     frame_buffer_pipeline_bridge_s1_arbiterlock2,
                                                     frame_buffer_pipeline_bridge_s1_burstcount,
                                                     frame_buffer_pipeline_bridge_s1_byteenable,
                                                     frame_buffer_pipeline_bridge_s1_chipselect,
                                                     frame_buffer_pipeline_bridge_s1_debugaccess,
                                                     frame_buffer_pipeline_bridge_s1_endofpacket_from_sa,
                                                     frame_buffer_pipeline_bridge_s1_nativeaddress,
                                                     frame_buffer_pipeline_bridge_s1_read,
                                                     frame_buffer_pipeline_bridge_s1_readdata_from_sa,
                                                     frame_buffer_pipeline_bridge_s1_reset_n,
                                                     frame_buffer_pipeline_bridge_s1_waitrequest_from_sa,
                                                     frame_buffer_pipeline_bridge_s1_write,
                                                     frame_buffer_pipeline_bridge_s1_writedata,
                                                     lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1,
                                                     lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1,
                                                     lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1,
                                                     lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                                     lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1,
                                                     pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1,
                                                     pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1,
                                                     pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1,
                                                     pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                                     pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1
                                                  )
;

  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1;
  output           accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1;
  output           d1_frame_buffer_pipeline_bridge_s1_end_xfer;
  output  [ 22: 0] frame_buffer_pipeline_bridge_s1_address;
  output           frame_buffer_pipeline_bridge_s1_arbiterlock;
  output           frame_buffer_pipeline_bridge_s1_arbiterlock2;
  output           frame_buffer_pipeline_bridge_s1_burstcount;
  output  [  3: 0] frame_buffer_pipeline_bridge_s1_byteenable;
  output           frame_buffer_pipeline_bridge_s1_chipselect;
  output           frame_buffer_pipeline_bridge_s1_debugaccess;
  output           frame_buffer_pipeline_bridge_s1_endofpacket_from_sa;
  output  [ 22: 0] frame_buffer_pipeline_bridge_s1_nativeaddress;
  output           frame_buffer_pipeline_bridge_s1_read;
  output  [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata_from_sa;
  output           frame_buffer_pipeline_bridge_s1_reset_n;
  output           frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;
  output           frame_buffer_pipeline_bridge_s1_write;
  output  [ 31: 0] frame_buffer_pipeline_bridge_s1_writedata;
  output           lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1;
  output           lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1;
  output           lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1;
  output           lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  output           lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1;
  output           pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1;
  output           pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1;
  output           pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1;
  output           pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  output           pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave;
  input   [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable;
  input            accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write;
  input   [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata;
  input            clk;
  input            frame_buffer_pipeline_bridge_s1_endofpacket;
  input   [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata;
  input            frame_buffer_pipeline_bridge_s1_readdatavalid;
  input            frame_buffer_pipeline_bridge_s1_waitrequest;
  input   [ 31: 0] lcd_sgdma_m_read_address_to_slave;
  input            lcd_sgdma_m_read_latency_counter;
  input            lcd_sgdma_m_read_read;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_debugaccess;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_saved_grant_frame_buffer_pipeline_bridge_s1;
  reg              d1_frame_buffer_pipeline_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1;
  wire    [ 22: 0] frame_buffer_pipeline_bridge_s1_address;
  wire             frame_buffer_pipeline_bridge_s1_allgrants;
  wire             frame_buffer_pipeline_bridge_s1_allow_new_arb_cycle;
  wire             frame_buffer_pipeline_bridge_s1_any_bursting_master_saved_grant;
  wire             frame_buffer_pipeline_bridge_s1_any_continuerequest;
  reg     [  2: 0] frame_buffer_pipeline_bridge_s1_arb_addend;
  wire             frame_buffer_pipeline_bridge_s1_arb_counter_enable;
  reg     [  6: 0] frame_buffer_pipeline_bridge_s1_arb_share_counter;
  wire    [  6: 0] frame_buffer_pipeline_bridge_s1_arb_share_counter_next_value;
  wire    [  6: 0] frame_buffer_pipeline_bridge_s1_arb_share_set_values;
  wire    [  2: 0] frame_buffer_pipeline_bridge_s1_arb_winner;
  wire             frame_buffer_pipeline_bridge_s1_arbiterlock;
  wire             frame_buffer_pipeline_bridge_s1_arbiterlock2;
  wire             frame_buffer_pipeline_bridge_s1_arbitration_holdoff_internal;
  wire             frame_buffer_pipeline_bridge_s1_beginbursttransfer_internal;
  wire             frame_buffer_pipeline_bridge_s1_begins_xfer;
  wire             frame_buffer_pipeline_bridge_s1_burstcount;
  wire    [  3: 0] frame_buffer_pipeline_bridge_s1_byteenable;
  wire             frame_buffer_pipeline_bridge_s1_chipselect;
  wire    [  5: 0] frame_buffer_pipeline_bridge_s1_chosen_master_double_vector;
  wire    [  2: 0] frame_buffer_pipeline_bridge_s1_chosen_master_rot_left;
  wire             frame_buffer_pipeline_bridge_s1_debugaccess;
  wire             frame_buffer_pipeline_bridge_s1_end_xfer;
  wire             frame_buffer_pipeline_bridge_s1_endofpacket_from_sa;
  wire             frame_buffer_pipeline_bridge_s1_firsttransfer;
  wire    [  2: 0] frame_buffer_pipeline_bridge_s1_grant_vector;
  wire             frame_buffer_pipeline_bridge_s1_in_a_read_cycle;
  wire             frame_buffer_pipeline_bridge_s1_in_a_write_cycle;
  wire    [  2: 0] frame_buffer_pipeline_bridge_s1_master_qreq_vector;
  wire             frame_buffer_pipeline_bridge_s1_move_on_to_next_transaction;
  wire    [ 22: 0] frame_buffer_pipeline_bridge_s1_nativeaddress;
  wire             frame_buffer_pipeline_bridge_s1_non_bursting_master_requests;
  wire             frame_buffer_pipeline_bridge_s1_read;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata_from_sa;
  wire             frame_buffer_pipeline_bridge_s1_readdatavalid_from_sa;
  reg              frame_buffer_pipeline_bridge_s1_reg_firsttransfer;
  wire             frame_buffer_pipeline_bridge_s1_reset_n;
  reg     [  2: 0] frame_buffer_pipeline_bridge_s1_saved_chosen_master_vector;
  reg              frame_buffer_pipeline_bridge_s1_slavearbiterlockenable;
  wire             frame_buffer_pipeline_bridge_s1_slavearbiterlockenable2;
  wire             frame_buffer_pipeline_bridge_s1_unreg_firsttransfer;
  wire             frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;
  wire             frame_buffer_pipeline_bridge_s1_waits_for_read;
  wire             frame_buffer_pipeline_bridge_s1_waits_for_write;
  wire             frame_buffer_pipeline_bridge_s1_write;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_s1_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_slave_frame_buffer_pipeline_bridge_s1;
  reg              last_cycle_lcd_sgdma_m_read_granted_slave_frame_buffer_pipeline_bridge_s1;
  reg              last_cycle_pipeline_bridge_m1_granted_slave_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_arbiterlock;
  wire             lcd_sgdma_m_read_arbiterlock2;
  wire             lcd_sgdma_m_read_continuerequest;
  wire             lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_rdv_fifo_output_from_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  wire             lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_saved_grant_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_rdv_fifo_output_from_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  wire             pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_saved_grant_frame_buffer_pipeline_bridge_s1;
  wire    [ 31: 0] shifted_address_to_frame_buffer_pipeline_bridge_s1_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1;
  wire    [ 31: 0] shifted_address_to_frame_buffer_pipeline_bridge_s1_from_lcd_sgdma_m_read;
  wire    [ 26: 0] shifted_address_to_frame_buffer_pipeline_bridge_s1_from_pipeline_bridge_m1;
  wire             wait_for_frame_buffer_pipeline_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~frame_buffer_pipeline_bridge_s1_end_xfer;
    end


  assign frame_buffer_pipeline_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1 | lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1 | pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1));
  //assign frame_buffer_pipeline_bridge_s1_readdatavalid_from_sa = frame_buffer_pipeline_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_readdatavalid_from_sa = frame_buffer_pipeline_bridge_s1_readdatavalid;

  //assign frame_buffer_pipeline_bridge_s1_readdata_from_sa = frame_buffer_pipeline_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_readdata_from_sa = frame_buffer_pipeline_bridge_s1_readdata;

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1 = (({accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave[31 : 25] , 25'b0} == 32'h0) & (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write)) & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write;
  //assign frame_buffer_pipeline_bridge_s1_waitrequest_from_sa = frame_buffer_pipeline_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_waitrequest_from_sa = frame_buffer_pipeline_bridge_s1_waitrequest;

  //frame_buffer_pipeline_bridge_s1_arb_share_counter set values, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_arb_share_set_values = (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1)? 100 :
    (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1)? 100 :
    (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1)? 100 :
    (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1)? 100 :
    1;

  //frame_buffer_pipeline_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_non_bursting_master_requests = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1 |
    lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1 |
    pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1 |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1 |
    lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1 |
    pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1 |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1 |
    lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1 |
    pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1 |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1 |
    lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1 |
    pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1;

  //frame_buffer_pipeline_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_any_bursting_master_saved_grant = 0;

  //frame_buffer_pipeline_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_arb_share_counter_next_value = frame_buffer_pipeline_bridge_s1_firsttransfer ? (frame_buffer_pipeline_bridge_s1_arb_share_set_values - 1) : |frame_buffer_pipeline_bridge_s1_arb_share_counter ? (frame_buffer_pipeline_bridge_s1_arb_share_counter - 1) : 0;

  //frame_buffer_pipeline_bridge_s1_allgrants all slave grants, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_allgrants = (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector) |
    (|frame_buffer_pipeline_bridge_s1_grant_vector);

  //frame_buffer_pipeline_bridge_s1_end_xfer assignment, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_end_xfer = ~(frame_buffer_pipeline_bridge_s1_waits_for_read | frame_buffer_pipeline_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_end_xfer & (~frame_buffer_pipeline_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //frame_buffer_pipeline_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1 & frame_buffer_pipeline_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1 & ~frame_buffer_pipeline_bridge_s1_non_bursting_master_requests);

  //frame_buffer_pipeline_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_s1_arb_share_counter <= 0;
      else if (frame_buffer_pipeline_bridge_s1_arb_counter_enable)
          frame_buffer_pipeline_bridge_s1_arb_share_counter <= frame_buffer_pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //frame_buffer_pipeline_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|frame_buffer_pipeline_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1) | (end_xfer_arb_share_counter_term_frame_buffer_pipeline_bridge_s1 & ~frame_buffer_pipeline_bridge_s1_non_bursting_master_requests))
          frame_buffer_pipeline_bridge_s1_slavearbiterlockenable <= |frame_buffer_pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 frame_buffer_pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock = frame_buffer_pipeline_bridge_s1_slavearbiterlockenable & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest;

  //frame_buffer_pipeline_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_slavearbiterlockenable2 = |frame_buffer_pipeline_bridge_s1_arb_share_counter_next_value;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 frame_buffer_pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock2 = frame_buffer_pipeline_bridge_s1_slavearbiterlockenable2 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest;

  //lcd_sgdma/m_read frame_buffer_pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign lcd_sgdma_m_read_arbiterlock = frame_buffer_pipeline_bridge_s1_slavearbiterlockenable & lcd_sgdma_m_read_continuerequest;

  //lcd_sgdma/m_read frame_buffer_pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign lcd_sgdma_m_read_arbiterlock2 = frame_buffer_pipeline_bridge_s1_slavearbiterlockenable2 & lcd_sgdma_m_read_continuerequest;

  //lcd_sgdma/m_read granted frame_buffer_pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_lcd_sgdma_m_read_granted_slave_frame_buffer_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_lcd_sgdma_m_read_granted_slave_frame_buffer_pipeline_bridge_s1 <= lcd_sgdma_m_read_saved_grant_frame_buffer_pipeline_bridge_s1 ? 1 : (frame_buffer_pipeline_bridge_s1_arbitration_holdoff_internal | ~lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1) ? 0 : last_cycle_lcd_sgdma_m_read_granted_slave_frame_buffer_pipeline_bridge_s1;
    end


  //lcd_sgdma_m_read_continuerequest continued request, which is an e_mux
  assign lcd_sgdma_m_read_continuerequest = (last_cycle_lcd_sgdma_m_read_granted_slave_frame_buffer_pipeline_bridge_s1 & lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1) |
    (last_cycle_lcd_sgdma_m_read_granted_slave_frame_buffer_pipeline_bridge_s1 & lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1);

  //frame_buffer_pipeline_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_any_continuerequest = lcd_sgdma_m_read_continuerequest |
    pipeline_bridge_m1_continuerequest |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest |
    pipeline_bridge_m1_continuerequest |
    accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest |
    lcd_sgdma_m_read_continuerequest;

  //pipeline_bridge/m1 frame_buffer_pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = frame_buffer_pipeline_bridge_s1_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //pipeline_bridge/m1 frame_buffer_pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = frame_buffer_pipeline_bridge_s1_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //pipeline_bridge/m1 granted frame_buffer_pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_pipeline_bridge_m1_granted_slave_frame_buffer_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_pipeline_bridge_m1_granted_slave_frame_buffer_pipeline_bridge_s1 <= pipeline_bridge_m1_saved_grant_frame_buffer_pipeline_bridge_s1 ? 1 : (frame_buffer_pipeline_bridge_s1_arbitration_holdoff_internal | ~pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1) ? 0 : last_cycle_pipeline_bridge_m1_granted_slave_frame_buffer_pipeline_bridge_s1;
    end


  //pipeline_bridge_m1_continuerequest continued request, which is an e_mux
  assign pipeline_bridge_m1_continuerequest = (last_cycle_pipeline_bridge_m1_granted_slave_frame_buffer_pipeline_bridge_s1 & pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1) |
    (last_cycle_pipeline_bridge_m1_granted_slave_frame_buffer_pipeline_bridge_s1 & pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1);

  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1 & ~(lcd_sgdma_m_read_arbiterlock | pipeline_bridge_m1_arbiterlock);
  //frame_buffer_pipeline_bridge_s1_writedata mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_writedata = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1)? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata :
    pipeline_bridge_m1_writedata;

  //assign frame_buffer_pipeline_bridge_s1_endofpacket_from_sa = frame_buffer_pipeline_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_endofpacket_from_sa = frame_buffer_pipeline_bridge_s1_endofpacket;

  assign lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1 = (({lcd_sgdma_m_read_address_to_slave[31 : 25] , 25'b0} == 32'h0) & (lcd_sgdma_m_read_read)) & lcd_sgdma_m_read_read;
  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 granted frame_buffer_pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_slave_frame_buffer_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_slave_frame_buffer_pipeline_bridge_s1 <= accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_saved_grant_frame_buffer_pipeline_bridge_s1 ? 1 : (frame_buffer_pipeline_bridge_s1_arbitration_holdoff_internal | ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1) ? 0 : last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_slave_frame_buffer_pipeline_bridge_s1;
    end


  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest continued request, which is an e_mux
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_continuerequest = (last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_slave_frame_buffer_pipeline_bridge_s1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1) |
    (last_cycle_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_slave_frame_buffer_pipeline_bridge_s1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1);

  assign lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1 = lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1 & ~((lcd_sgdma_m_read_read & ((lcd_sgdma_m_read_latency_counter != 0) | (1 < lcd_sgdma_m_read_latency_counter))) | accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock | pipeline_bridge_m1_arbiterlock);
  //unique name for frame_buffer_pipeline_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_move_on_to_next_transaction = frame_buffer_pipeline_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_lcd_sgdma_m_read_to_frame_buffer_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_lcd_sgdma_m_read_to_frame_buffer_pipeline_bridge_s1_module rdv_fifo_for_lcd_sgdma_m_read_to_frame_buffer_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1),
      .data_out             (lcd_sgdma_m_read_rdv_fifo_output_from_frame_buffer_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (lcd_sgdma_m_read_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1),
      .full                 (),
      .read                 (frame_buffer_pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~frame_buffer_pipeline_bridge_s1_waits_for_read)
    );

  assign lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register = ~lcd_sgdma_m_read_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1;
  //local readdatavalid lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1, which is an e_mux
  assign lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1 = (frame_buffer_pipeline_bridge_s1_readdatavalid_from_sa & lcd_sgdma_m_read_rdv_fifo_output_from_frame_buffer_pipeline_bridge_s1) & ~ lcd_sgdma_m_read_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1;

  assign pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1 = ({pipeline_bridge_m1_address_to_slave[26 : 25] , 25'b0} == 27'h0) & pipeline_bridge_m1_chipselect;
  assign pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1 = pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1 & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0) | (1 < pipeline_bridge_m1_latency_counter) | (|pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register))) | accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock | lcd_sgdma_m_read_arbiterlock);
  //rdv_fifo_for_pipeline_bridge_m1_to_frame_buffer_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pipeline_bridge_m1_to_frame_buffer_pipeline_bridge_s1_module rdv_fifo_for_pipeline_bridge_m1_to_frame_buffer_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1),
      .data_out             (pipeline_bridge_m1_rdv_fifo_output_from_frame_buffer_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (pipeline_bridge_m1_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1),
      .full                 (),
      .read                 (frame_buffer_pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~frame_buffer_pipeline_bridge_s1_waits_for_read)
    );

  assign pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register = ~pipeline_bridge_m1_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1;
  //local readdatavalid pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1 = (frame_buffer_pipeline_bridge_s1_readdatavalid_from_sa & pipeline_bridge_m1_rdv_fifo_output_from_frame_buffer_pipeline_bridge_s1) & ~ pipeline_bridge_m1_rdv_fifo_empty_frame_buffer_pipeline_bridge_s1;

  //allow new arb cycle for frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_allow_new_arb_cycle = ~accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock & ~lcd_sgdma_m_read_arbiterlock & ~pipeline_bridge_m1_arbiterlock;

  //pipeline_bridge/m1 assignment into master qualified-requests vector for frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_master_qreq_vector[0] = pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1;

  //pipeline_bridge/m1 grant frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_grant_vector[0];

  //pipeline_bridge/m1 saved-grant frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_arb_winner[0] && pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1;

  //lcd_sgdma/m_read assignment into master qualified-requests vector for frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_master_qreq_vector[1] = lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1;

  //lcd_sgdma/m_read grant frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_grant_vector[1];

  //lcd_sgdma/m_read saved-grant frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign lcd_sgdma_m_read_saved_grant_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_arb_winner[1] && lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 assignment into master qualified-requests vector for frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_master_qreq_vector[2] = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1;

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 grant frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_grant_vector[2];

  //accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance/accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 saved-grant frame_buffer_pipeline_bridge/s1, which is an e_assign
  assign accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_saved_grant_frame_buffer_pipeline_bridge_s1 = frame_buffer_pipeline_bridge_s1_arb_winner[2] && accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1;

  //frame_buffer_pipeline_bridge/s1 chosen-master double-vector, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_chosen_master_double_vector = {frame_buffer_pipeline_bridge_s1_master_qreq_vector, frame_buffer_pipeline_bridge_s1_master_qreq_vector} & ({~frame_buffer_pipeline_bridge_s1_master_qreq_vector, ~frame_buffer_pipeline_bridge_s1_master_qreq_vector} + frame_buffer_pipeline_bridge_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign frame_buffer_pipeline_bridge_s1_arb_winner = (frame_buffer_pipeline_bridge_s1_allow_new_arb_cycle & | frame_buffer_pipeline_bridge_s1_grant_vector) ? frame_buffer_pipeline_bridge_s1_grant_vector : frame_buffer_pipeline_bridge_s1_saved_chosen_master_vector;

  //saved frame_buffer_pipeline_bridge_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_s1_saved_chosen_master_vector <= 0;
      else if (frame_buffer_pipeline_bridge_s1_allow_new_arb_cycle)
          frame_buffer_pipeline_bridge_s1_saved_chosen_master_vector <= |frame_buffer_pipeline_bridge_s1_grant_vector ? frame_buffer_pipeline_bridge_s1_grant_vector : frame_buffer_pipeline_bridge_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign frame_buffer_pipeline_bridge_s1_grant_vector = {(frame_buffer_pipeline_bridge_s1_chosen_master_double_vector[2] | frame_buffer_pipeline_bridge_s1_chosen_master_double_vector[5]),
    (frame_buffer_pipeline_bridge_s1_chosen_master_double_vector[1] | frame_buffer_pipeline_bridge_s1_chosen_master_double_vector[4]),
    (frame_buffer_pipeline_bridge_s1_chosen_master_double_vector[0] | frame_buffer_pipeline_bridge_s1_chosen_master_double_vector[3])};

  //frame_buffer_pipeline_bridge/s1 chosen master rotated left, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_chosen_master_rot_left = (frame_buffer_pipeline_bridge_s1_arb_winner << 1) ? (frame_buffer_pipeline_bridge_s1_arb_winner << 1) : 1;

  //frame_buffer_pipeline_bridge/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_s1_arb_addend <= 1;
      else if (|frame_buffer_pipeline_bridge_s1_grant_vector)
          frame_buffer_pipeline_bridge_s1_arb_addend <= frame_buffer_pipeline_bridge_s1_end_xfer? frame_buffer_pipeline_bridge_s1_chosen_master_rot_left : frame_buffer_pipeline_bridge_s1_grant_vector;
    end


  //frame_buffer_pipeline_bridge_s1_reset_n assignment, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_reset_n = reset_n;

  assign frame_buffer_pipeline_bridge_s1_chipselect = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1 | lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1 | pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1;
  //frame_buffer_pipeline_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_firsttransfer = frame_buffer_pipeline_bridge_s1_begins_xfer ? frame_buffer_pipeline_bridge_s1_unreg_firsttransfer : frame_buffer_pipeline_bridge_s1_reg_firsttransfer;

  //frame_buffer_pipeline_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_unreg_firsttransfer = ~(frame_buffer_pipeline_bridge_s1_slavearbiterlockenable & frame_buffer_pipeline_bridge_s1_any_continuerequest);

  //frame_buffer_pipeline_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (frame_buffer_pipeline_bridge_s1_begins_xfer)
          frame_buffer_pipeline_bridge_s1_reg_firsttransfer <= frame_buffer_pipeline_bridge_s1_unreg_firsttransfer;
    end


  //frame_buffer_pipeline_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_beginbursttransfer_internal = frame_buffer_pipeline_bridge_s1_begins_xfer;

  //frame_buffer_pipeline_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_arbitration_holdoff_internal = frame_buffer_pipeline_bridge_s1_begins_xfer & frame_buffer_pipeline_bridge_s1_firsttransfer;

  //frame_buffer_pipeline_bridge_s1_read assignment, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_read = (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1 & lcd_sgdma_m_read_read) | (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect));

  //frame_buffer_pipeline_bridge_s1_write assignment, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_write = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write) | (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect));

  assign shifted_address_to_frame_buffer_pipeline_bridge_s1_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 = accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave;
  //frame_buffer_pipeline_bridge_s1_address mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_address = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1)? (shifted_address_to_frame_buffer_pipeline_bridge_s1_from_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1 >> 2) :
    (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1)? (shifted_address_to_frame_buffer_pipeline_bridge_s1_from_lcd_sgdma_m_read >> 2) :
    (shifted_address_to_frame_buffer_pipeline_bridge_s1_from_pipeline_bridge_m1 >> 2);

  assign shifted_address_to_frame_buffer_pipeline_bridge_s1_from_lcd_sgdma_m_read = lcd_sgdma_m_read_address_to_slave;
  assign shifted_address_to_frame_buffer_pipeline_bridge_s1_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //slaveid frame_buffer_pipeline_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_nativeaddress = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1)? (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave >> 2) :
    (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1)? (lcd_sgdma_m_read_address_to_slave >> 2) :
    (pipeline_bridge_m1_address_to_slave >> 2);

  //d1_frame_buffer_pipeline_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_frame_buffer_pipeline_bridge_s1_end_xfer <= 1;
      else 
        d1_frame_buffer_pipeline_bridge_s1_end_xfer <= frame_buffer_pipeline_bridge_s1_end_xfer;
    end


  //frame_buffer_pipeline_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_waits_for_read = frame_buffer_pipeline_bridge_s1_in_a_read_cycle & frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;

  //frame_buffer_pipeline_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_in_a_read_cycle = (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1 & lcd_sgdma_m_read_read) | (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect));

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = frame_buffer_pipeline_bridge_s1_in_a_read_cycle;

  //frame_buffer_pipeline_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_waits_for_write = frame_buffer_pipeline_bridge_s1_in_a_write_cycle & frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;

  //frame_buffer_pipeline_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign frame_buffer_pipeline_bridge_s1_in_a_write_cycle = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1 & accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write) | (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect));

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = frame_buffer_pipeline_bridge_s1_in_a_write_cycle;

  assign wait_for_frame_buffer_pipeline_bridge_s1_counter = 0;
  //frame_buffer_pipeline_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_byteenable = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1)? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable :
    (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1)? pipeline_bridge_m1_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_burstcount = (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1)? pipeline_bridge_m1_burstcount :
    1;

  //frame_buffer_pipeline_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_arbiterlock = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock)? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock :
    (lcd_sgdma_m_read_arbiterlock)? lcd_sgdma_m_read_arbiterlock :
    pipeline_bridge_m1_arbiterlock;

  //frame_buffer_pipeline_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_arbiterlock2 = (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock2)? accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbiterlock2 :
    (lcd_sgdma_m_read_arbiterlock2)? lcd_sgdma_m_read_arbiterlock2 :
    pipeline_bridge_m1_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_s1_debugaccess = (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1)? pipeline_bridge_m1_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //frame_buffer_pipeline_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1 && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave frame_buffer_pipeline_bridge/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1 + lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1 + pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_saved_grant_frame_buffer_pipeline_bridge_s1 + lcd_sgdma_m_read_saved_grant_frame_buffer_pipeline_bridge_s1 + pipeline_bridge_m1_saved_grant_frame_buffer_pipeline_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module frame_buffer_pipeline_bridge_m1_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer,
                                                     ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa,
                                                     ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa,
                                                     ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa,
                                                     frame_buffer_pipeline_bridge_m1_address,
                                                     frame_buffer_pipeline_bridge_m1_burstcount,
                                                     frame_buffer_pipeline_bridge_m1_byteenable,
                                                     frame_buffer_pipeline_bridge_m1_chipselect,
                                                     frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1,
                                                     frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1,
                                                     frame_buffer_pipeline_bridge_m1_read,
                                                     frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1,
                                                     frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register,
                                                     frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1,
                                                     frame_buffer_pipeline_bridge_m1_write,
                                                     frame_buffer_pipeline_bridge_m1_writedata,
                                                     reset_n,

                                                    // outputs:
                                                     frame_buffer_pipeline_bridge_m1_address_to_slave,
                                                     frame_buffer_pipeline_bridge_m1_endofpacket,
                                                     frame_buffer_pipeline_bridge_m1_latency_counter,
                                                     frame_buffer_pipeline_bridge_m1_readdata,
                                                     frame_buffer_pipeline_bridge_m1_readdatavalid,
                                                     frame_buffer_pipeline_bridge_m1_waitrequest
                                                  )
;

  output  [ 24: 0] frame_buffer_pipeline_bridge_m1_address_to_slave;
  output           frame_buffer_pipeline_bridge_m1_endofpacket;
  output           frame_buffer_pipeline_bridge_m1_latency_counter;
  output  [ 31: 0] frame_buffer_pipeline_bridge_m1_readdata;
  output           frame_buffer_pipeline_bridge_m1_readdatavalid;
  output           frame_buffer_pipeline_bridge_m1_waitrequest;
  input            clk;
  input            d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer;
  input            ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa;
  input   [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa;
  input            ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa;
  input   [ 24: 0] frame_buffer_pipeline_bridge_m1_address;
  input            frame_buffer_pipeline_bridge_m1_burstcount;
  input   [  3: 0] frame_buffer_pipeline_bridge_m1_byteenable;
  input            frame_buffer_pipeline_bridge_m1_chipselect;
  input            frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1;
  input            frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1;
  input            frame_buffer_pipeline_bridge_m1_read;
  input            frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1;
  input            frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register;
  input            frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1;
  input            frame_buffer_pipeline_bridge_m1_write;
  input   [ 31: 0] frame_buffer_pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] frame_buffer_pipeline_bridge_m1_address_last_time;
  wire    [ 24: 0] frame_buffer_pipeline_bridge_m1_address_to_slave;
  reg              frame_buffer_pipeline_bridge_m1_burstcount_last_time;
  reg     [  3: 0] frame_buffer_pipeline_bridge_m1_byteenable_last_time;
  reg              frame_buffer_pipeline_bridge_m1_chipselect_last_time;
  wire             frame_buffer_pipeline_bridge_m1_endofpacket;
  wire             frame_buffer_pipeline_bridge_m1_latency_counter;
  reg              frame_buffer_pipeline_bridge_m1_read_last_time;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_m1_readdata;
  wire             frame_buffer_pipeline_bridge_m1_readdatavalid;
  wire             frame_buffer_pipeline_bridge_m1_run;
  wire             frame_buffer_pipeline_bridge_m1_waitrequest;
  reg              frame_buffer_pipeline_bridge_m1_write_last_time;
  reg     [ 31: 0] frame_buffer_pipeline_bridge_m1_writedata_last_time;
  wire             pre_flush_frame_buffer_pipeline_bridge_m1_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1 | ~frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1) & ((~frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1 | ~frame_buffer_pipeline_bridge_m1_chipselect | (1 & ~ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa & frame_buffer_pipeline_bridge_m1_chipselect))) & ((~frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1 | ~frame_buffer_pipeline_bridge_m1_chipselect | (1 & ~ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa & frame_buffer_pipeline_bridge_m1_chipselect)));

  //cascaded wait assignment, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign frame_buffer_pipeline_bridge_m1_address_to_slave = frame_buffer_pipeline_bridge_m1_address[24 : 0];

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_frame_buffer_pipeline_bridge_m1_readdatavalid = frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign frame_buffer_pipeline_bridge_m1_readdatavalid = 0 |
    pre_flush_frame_buffer_pipeline_bridge_m1_readdatavalid;

  //frame_buffer_pipeline_bridge/m1 readdata mux, which is an e_mux
  assign frame_buffer_pipeline_bridge_m1_readdata = ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_waitrequest = ~frame_buffer_pipeline_bridge_m1_run;

  //latent max counter, which is an e_assign
  assign frame_buffer_pipeline_bridge_m1_latency_counter = 0;

  //mux frame_buffer_pipeline_bridge_m1_endofpacket, which is an e_mux
  assign frame_buffer_pipeline_bridge_m1_endofpacket = ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //frame_buffer_pipeline_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_address_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_address_last_time <= frame_buffer_pipeline_bridge_m1_address;
    end


  //frame_buffer_pipeline_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= frame_buffer_pipeline_bridge_m1_waitrequest & frame_buffer_pipeline_bridge_m1_chipselect;
    end


  //frame_buffer_pipeline_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_address != frame_buffer_pipeline_bridge_m1_address_last_time))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //frame_buffer_pipeline_bridge_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_chipselect_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_chipselect_last_time <= frame_buffer_pipeline_bridge_m1_chipselect;
    end


  //frame_buffer_pipeline_bridge_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_chipselect != frame_buffer_pipeline_bridge_m1_chipselect_last_time))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //frame_buffer_pipeline_bridge_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_burstcount_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_burstcount_last_time <= frame_buffer_pipeline_bridge_m1_burstcount;
    end


  //frame_buffer_pipeline_bridge_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_burstcount != frame_buffer_pipeline_bridge_m1_burstcount_last_time))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //frame_buffer_pipeline_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_byteenable_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_byteenable_last_time <= frame_buffer_pipeline_bridge_m1_byteenable;
    end


  //frame_buffer_pipeline_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_byteenable != frame_buffer_pipeline_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //frame_buffer_pipeline_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_read_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_read_last_time <= frame_buffer_pipeline_bridge_m1_read;
    end


  //frame_buffer_pipeline_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_read != frame_buffer_pipeline_bridge_m1_read_last_time))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //frame_buffer_pipeline_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_write_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_write_last_time <= frame_buffer_pipeline_bridge_m1_write;
    end


  //frame_buffer_pipeline_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_write != frame_buffer_pipeline_bridge_m1_write_last_time))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //frame_buffer_pipeline_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          frame_buffer_pipeline_bridge_m1_writedata_last_time <= 0;
      else 
        frame_buffer_pipeline_bridge_m1_writedata_last_time <= frame_buffer_pipeline_bridge_m1_writedata;
    end


  //frame_buffer_pipeline_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (frame_buffer_pipeline_bridge_m1_writedata != frame_buffer_pipeline_bridge_m1_writedata_last_time) & (frame_buffer_pipeline_bridge_m1_write & frame_buffer_pipeline_bridge_m1_chipselect))
        begin
          $write("%0d ns: frame_buffer_pipeline_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module frame_buffer_pipeline_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 clock_crossing_bridge_m1_address_to_slave,
                                                 clock_crossing_bridge_m1_latency_counter,
                                                 clock_crossing_bridge_m1_nativeaddress,
                                                 clock_crossing_bridge_m1_read,
                                                 clock_crossing_bridge_m1_write,
                                                 clock_crossing_bridge_m1_writedata,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
                                                 clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata
                                              )
;

  output           clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  output           clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  output           clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave;
  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg              jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire             jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire             jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave = ({clock_crossing_bridge_m1_address_to_slave[10 : 3] , 3'b0} == 11'h580) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave = clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave = clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave & clock_crossing_bridge_m1_read & ~jtag_uart_avalon_jtag_slave_waits_for_read;

  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave = clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;

  //clock_crossing_bridge/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave = clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave & clock_crossing_bridge_m1_read);

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave & clock_crossing_bridge_m1_write);

  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_data_format_adapter_in_arbitrator (
                                               // inputs:
                                                clk,
                                                lcd_data_format_adapter_in_ready,
                                                lcd_pixel_converter_out_data,
                                                lcd_pixel_converter_out_empty,
                                                lcd_pixel_converter_out_endofpacket,
                                                lcd_pixel_converter_out_startofpacket,
                                                lcd_pixel_converter_out_valid,
                                                reset_n,

                                               // outputs:
                                                lcd_data_format_adapter_in_data,
                                                lcd_data_format_adapter_in_empty,
                                                lcd_data_format_adapter_in_endofpacket,
                                                lcd_data_format_adapter_in_ready_from_sa,
                                                lcd_data_format_adapter_in_reset_n,
                                                lcd_data_format_adapter_in_startofpacket,
                                                lcd_data_format_adapter_in_valid
                                             )
;

  output  [ 23: 0] lcd_data_format_adapter_in_data;
  output  [  1: 0] lcd_data_format_adapter_in_empty;
  output           lcd_data_format_adapter_in_endofpacket;
  output           lcd_data_format_adapter_in_ready_from_sa;
  output           lcd_data_format_adapter_in_reset_n;
  output           lcd_data_format_adapter_in_startofpacket;
  output           lcd_data_format_adapter_in_valid;
  input            clk;
  input            lcd_data_format_adapter_in_ready;
  input   [ 23: 0] lcd_pixel_converter_out_data;
  input   [  1: 0] lcd_pixel_converter_out_empty;
  input            lcd_pixel_converter_out_endofpacket;
  input            lcd_pixel_converter_out_startofpacket;
  input            lcd_pixel_converter_out_valid;
  input            reset_n;

  wire    [ 23: 0] lcd_data_format_adapter_in_data;
  wire    [  1: 0] lcd_data_format_adapter_in_empty;
  wire             lcd_data_format_adapter_in_endofpacket;
  wire             lcd_data_format_adapter_in_ready_from_sa;
  wire             lcd_data_format_adapter_in_reset_n;
  wire             lcd_data_format_adapter_in_startofpacket;
  wire             lcd_data_format_adapter_in_valid;
  //mux lcd_data_format_adapter_in_data, which is an e_mux
  assign lcd_data_format_adapter_in_data = lcd_pixel_converter_out_data;

  //mux lcd_data_format_adapter_in_empty, which is an e_mux
  assign lcd_data_format_adapter_in_empty = lcd_pixel_converter_out_empty;

  //mux lcd_data_format_adapter_in_endofpacket, which is an e_mux
  assign lcd_data_format_adapter_in_endofpacket = lcd_pixel_converter_out_endofpacket;

  //assign lcd_data_format_adapter_in_ready_from_sa = lcd_data_format_adapter_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_data_format_adapter_in_ready_from_sa = lcd_data_format_adapter_in_ready;

  //mux lcd_data_format_adapter_in_startofpacket, which is an e_mux
  assign lcd_data_format_adapter_in_startofpacket = lcd_pixel_converter_out_startofpacket;

  //mux lcd_data_format_adapter_in_valid, which is an e_mux
  assign lcd_data_format_adapter_in_valid = lcd_pixel_converter_out_valid;

  //lcd_data_format_adapter_in_reset_n assignment, which is an e_assign
  assign lcd_data_format_adapter_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_data_format_adapter_out_arbitrator (
                                                // inputs:
                                                 clk,
                                                 lcd_data_format_adapter_out_data,
                                                 lcd_data_format_adapter_out_endofpacket,
                                                 lcd_data_format_adapter_out_startofpacket,
                                                 lcd_data_format_adapter_out_valid,
                                                 lcd_ta_formatter_to_fifo_in_ready_from_sa,
                                                 reset_n,

                                                // outputs:
                                                 lcd_data_format_adapter_out_ready
                                              )
;

  output           lcd_data_format_adapter_out_ready;
  input            clk;
  input   [  7: 0] lcd_data_format_adapter_out_data;
  input            lcd_data_format_adapter_out_endofpacket;
  input            lcd_data_format_adapter_out_startofpacket;
  input            lcd_data_format_adapter_out_valid;
  input            lcd_ta_formatter_to_fifo_in_ready_from_sa;
  input            reset_n;

  wire             lcd_data_format_adapter_out_ready;
  //mux lcd_data_format_adapter_out_ready, which is an e_mux
  assign lcd_data_format_adapter_out_ready = lcd_ta_formatter_to_fifo_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_data_format_adapter_1_in_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  lcd_data_format_adapter_1_in_ready,
                                                  lcd_ta_fifo_to_sequencer_out_data,
                                                  lcd_ta_fifo_to_sequencer_out_endofpacket,
                                                  lcd_ta_fifo_to_sequencer_out_startofpacket,
                                                  lcd_ta_fifo_to_sequencer_out_valid,
                                                  reset_n,

                                                 // outputs:
                                                  lcd_data_format_adapter_1_in_data,
                                                  lcd_data_format_adapter_1_in_endofpacket,
                                                  lcd_data_format_adapter_1_in_ready_from_sa,
                                                  lcd_data_format_adapter_1_in_reset_n,
                                                  lcd_data_format_adapter_1_in_startofpacket,
                                                  lcd_data_format_adapter_1_in_valid
                                               )
;

  output  [  7: 0] lcd_data_format_adapter_1_in_data;
  output           lcd_data_format_adapter_1_in_endofpacket;
  output           lcd_data_format_adapter_1_in_ready_from_sa;
  output           lcd_data_format_adapter_1_in_reset_n;
  output           lcd_data_format_adapter_1_in_startofpacket;
  output           lcd_data_format_adapter_1_in_valid;
  input            clk;
  input            lcd_data_format_adapter_1_in_ready;
  input   [  7: 0] lcd_ta_fifo_to_sequencer_out_data;
  input            lcd_ta_fifo_to_sequencer_out_endofpacket;
  input            lcd_ta_fifo_to_sequencer_out_startofpacket;
  input            lcd_ta_fifo_to_sequencer_out_valid;
  input            reset_n;

  wire    [  7: 0] lcd_data_format_adapter_1_in_data;
  wire             lcd_data_format_adapter_1_in_endofpacket;
  wire             lcd_data_format_adapter_1_in_ready_from_sa;
  wire             lcd_data_format_adapter_1_in_reset_n;
  wire             lcd_data_format_adapter_1_in_startofpacket;
  wire             lcd_data_format_adapter_1_in_valid;
  //mux lcd_data_format_adapter_1_in_data, which is an e_mux
  assign lcd_data_format_adapter_1_in_data = lcd_ta_fifo_to_sequencer_out_data;

  //mux lcd_data_format_adapter_1_in_endofpacket, which is an e_mux
  assign lcd_data_format_adapter_1_in_endofpacket = lcd_ta_fifo_to_sequencer_out_endofpacket;

  //assign lcd_data_format_adapter_1_in_ready_from_sa = lcd_data_format_adapter_1_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_data_format_adapter_1_in_ready_from_sa = lcd_data_format_adapter_1_in_ready;

  //mux lcd_data_format_adapter_1_in_startofpacket, which is an e_mux
  assign lcd_data_format_adapter_1_in_startofpacket = lcd_ta_fifo_to_sequencer_out_startofpacket;

  //mux lcd_data_format_adapter_1_in_valid, which is an e_mux
  assign lcd_data_format_adapter_1_in_valid = lcd_ta_fifo_to_sequencer_out_valid;

  //lcd_data_format_adapter_1_in_reset_n assignment, which is an e_assign
  assign lcd_data_format_adapter_1_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_data_format_adapter_1_out_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   lcd_data_format_adapter_1_out_data,
                                                   lcd_data_format_adapter_1_out_empty,
                                                   lcd_data_format_adapter_1_out_endofpacket,
                                                   lcd_data_format_adapter_1_out_startofpacket,
                                                   lcd_data_format_adapter_1_out_valid,
                                                   lcd_video_sequencer_in_ready_from_sa,
                                                   reset_n,

                                                  // outputs:
                                                   lcd_data_format_adapter_1_out_ready
                                                )
;

  output           lcd_data_format_adapter_1_out_ready;
  input            clk;
  input   [  7: 0] lcd_data_format_adapter_1_out_data;
  input            lcd_data_format_adapter_1_out_empty;
  input            lcd_data_format_adapter_1_out_endofpacket;
  input            lcd_data_format_adapter_1_out_startofpacket;
  input            lcd_data_format_adapter_1_out_valid;
  input            lcd_video_sequencer_in_ready_from_sa;
  input            reset_n;

  wire             lcd_data_format_adapter_1_out_ready;
  //mux lcd_data_format_adapter_1_out_ready, which is an e_mux
  assign lcd_data_format_adapter_1_out_ready = lcd_video_sequencer_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_i2c_cs_s1_arbitrator (
                                  // inputs:
                                   clk,
                                   clock_crossing_bridge_m1_address_to_slave,
                                   clock_crossing_bridge_m1_latency_counter,
                                   clock_crossing_bridge_m1_nativeaddress,
                                   clock_crossing_bridge_m1_read,
                                   clock_crossing_bridge_m1_write,
                                   clock_crossing_bridge_m1_writedata,
                                   lcd_i2c_cs_s1_readdata,
                                   reset_n,

                                  // outputs:
                                   clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1,
                                   clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1,
                                   clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1,
                                   clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1,
                                   d1_lcd_i2c_cs_s1_end_xfer,
                                   lcd_i2c_cs_s1_address,
                                   lcd_i2c_cs_s1_chipselect,
                                   lcd_i2c_cs_s1_readdata_from_sa,
                                   lcd_i2c_cs_s1_reset_n,
                                   lcd_i2c_cs_s1_write_n,
                                   lcd_i2c_cs_s1_writedata
                                )
;

  output           clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1;
  output           clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1;
  output           clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1;
  output           clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1;
  output           d1_lcd_i2c_cs_s1_end_xfer;
  output  [  1: 0] lcd_i2c_cs_s1_address;
  output           lcd_i2c_cs_s1_chipselect;
  output  [ 31: 0] lcd_i2c_cs_s1_readdata_from_sa;
  output           lcd_i2c_cs_s1_reset_n;
  output           lcd_i2c_cs_s1_write_n;
  output  [ 31: 0] lcd_i2c_cs_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] lcd_i2c_cs_s1_readdata;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_saved_grant_lcd_i2c_cs_s1;
  reg              d1_lcd_i2c_cs_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_lcd_i2c_cs_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] lcd_i2c_cs_s1_address;
  wire             lcd_i2c_cs_s1_allgrants;
  wire             lcd_i2c_cs_s1_allow_new_arb_cycle;
  wire             lcd_i2c_cs_s1_any_bursting_master_saved_grant;
  wire             lcd_i2c_cs_s1_any_continuerequest;
  wire             lcd_i2c_cs_s1_arb_counter_enable;
  reg              lcd_i2c_cs_s1_arb_share_counter;
  wire             lcd_i2c_cs_s1_arb_share_counter_next_value;
  wire             lcd_i2c_cs_s1_arb_share_set_values;
  wire             lcd_i2c_cs_s1_beginbursttransfer_internal;
  wire             lcd_i2c_cs_s1_begins_xfer;
  wire             lcd_i2c_cs_s1_chipselect;
  wire             lcd_i2c_cs_s1_end_xfer;
  wire             lcd_i2c_cs_s1_firsttransfer;
  wire             lcd_i2c_cs_s1_grant_vector;
  wire             lcd_i2c_cs_s1_in_a_read_cycle;
  wire             lcd_i2c_cs_s1_in_a_write_cycle;
  wire             lcd_i2c_cs_s1_master_qreq_vector;
  wire             lcd_i2c_cs_s1_non_bursting_master_requests;
  wire    [ 31: 0] lcd_i2c_cs_s1_readdata_from_sa;
  reg              lcd_i2c_cs_s1_reg_firsttransfer;
  wire             lcd_i2c_cs_s1_reset_n;
  reg              lcd_i2c_cs_s1_slavearbiterlockenable;
  wire             lcd_i2c_cs_s1_slavearbiterlockenable2;
  wire             lcd_i2c_cs_s1_unreg_firsttransfer;
  wire             lcd_i2c_cs_s1_waits_for_read;
  wire             lcd_i2c_cs_s1_waits_for_write;
  wire             lcd_i2c_cs_s1_write_n;
  wire    [ 31: 0] lcd_i2c_cs_s1_writedata;
  wire             wait_for_lcd_i2c_cs_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~lcd_i2c_cs_s1_end_xfer;
    end


  assign lcd_i2c_cs_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1));
  //assign lcd_i2c_cs_s1_readdata_from_sa = lcd_i2c_cs_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_i2c_cs_s1_readdata_from_sa = lcd_i2c_cs_s1_readdata;

  assign clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h380) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //lcd_i2c_cs_s1_arb_share_counter set values, which is an e_mux
  assign lcd_i2c_cs_s1_arb_share_set_values = 1;

  //lcd_i2c_cs_s1_non_bursting_master_requests mux, which is an e_mux
  assign lcd_i2c_cs_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1;

  //lcd_i2c_cs_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign lcd_i2c_cs_s1_any_bursting_master_saved_grant = 0;

  //lcd_i2c_cs_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign lcd_i2c_cs_s1_arb_share_counter_next_value = lcd_i2c_cs_s1_firsttransfer ? (lcd_i2c_cs_s1_arb_share_set_values - 1) : |lcd_i2c_cs_s1_arb_share_counter ? (lcd_i2c_cs_s1_arb_share_counter - 1) : 0;

  //lcd_i2c_cs_s1_allgrants all slave grants, which is an e_mux
  assign lcd_i2c_cs_s1_allgrants = |lcd_i2c_cs_s1_grant_vector;

  //lcd_i2c_cs_s1_end_xfer assignment, which is an e_assign
  assign lcd_i2c_cs_s1_end_xfer = ~(lcd_i2c_cs_s1_waits_for_read | lcd_i2c_cs_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_lcd_i2c_cs_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_lcd_i2c_cs_s1 = lcd_i2c_cs_s1_end_xfer & (~lcd_i2c_cs_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //lcd_i2c_cs_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign lcd_i2c_cs_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_lcd_i2c_cs_s1 & lcd_i2c_cs_s1_allgrants) | (end_xfer_arb_share_counter_term_lcd_i2c_cs_s1 & ~lcd_i2c_cs_s1_non_bursting_master_requests);

  //lcd_i2c_cs_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_cs_s1_arb_share_counter <= 0;
      else if (lcd_i2c_cs_s1_arb_counter_enable)
          lcd_i2c_cs_s1_arb_share_counter <= lcd_i2c_cs_s1_arb_share_counter_next_value;
    end


  //lcd_i2c_cs_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_cs_s1_slavearbiterlockenable <= 0;
      else if ((|lcd_i2c_cs_s1_master_qreq_vector & end_xfer_arb_share_counter_term_lcd_i2c_cs_s1) | (end_xfer_arb_share_counter_term_lcd_i2c_cs_s1 & ~lcd_i2c_cs_s1_non_bursting_master_requests))
          lcd_i2c_cs_s1_slavearbiterlockenable <= |lcd_i2c_cs_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 lcd_i2c_cs/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = lcd_i2c_cs_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //lcd_i2c_cs_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign lcd_i2c_cs_s1_slavearbiterlockenable2 = |lcd_i2c_cs_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 lcd_i2c_cs/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = lcd_i2c_cs_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //lcd_i2c_cs_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign lcd_i2c_cs_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1 = clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1 = clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1 & clock_crossing_bridge_m1_read & ~lcd_i2c_cs_s1_waits_for_read;

  //lcd_i2c_cs_s1_writedata mux, which is an e_mux
  assign lcd_i2c_cs_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1 = clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1;

  //clock_crossing_bridge/m1 saved-grant lcd_i2c_cs/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_lcd_i2c_cs_s1 = clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1;

  //allow new arb cycle for lcd_i2c_cs/s1, which is an e_assign
  assign lcd_i2c_cs_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign lcd_i2c_cs_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign lcd_i2c_cs_s1_master_qreq_vector = 1;

  //lcd_i2c_cs_s1_reset_n assignment, which is an e_assign
  assign lcd_i2c_cs_s1_reset_n = reset_n;

  assign lcd_i2c_cs_s1_chipselect = clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1;
  //lcd_i2c_cs_s1_firsttransfer first transaction, which is an e_assign
  assign lcd_i2c_cs_s1_firsttransfer = lcd_i2c_cs_s1_begins_xfer ? lcd_i2c_cs_s1_unreg_firsttransfer : lcd_i2c_cs_s1_reg_firsttransfer;

  //lcd_i2c_cs_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign lcd_i2c_cs_s1_unreg_firsttransfer = ~(lcd_i2c_cs_s1_slavearbiterlockenable & lcd_i2c_cs_s1_any_continuerequest);

  //lcd_i2c_cs_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_cs_s1_reg_firsttransfer <= 1'b1;
      else if (lcd_i2c_cs_s1_begins_xfer)
          lcd_i2c_cs_s1_reg_firsttransfer <= lcd_i2c_cs_s1_unreg_firsttransfer;
    end


  //lcd_i2c_cs_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign lcd_i2c_cs_s1_beginbursttransfer_internal = lcd_i2c_cs_s1_begins_xfer;

  //~lcd_i2c_cs_s1_write_n assignment, which is an e_mux
  assign lcd_i2c_cs_s1_write_n = ~(clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1 & clock_crossing_bridge_m1_write);

  //lcd_i2c_cs_s1_address mux, which is an e_mux
  assign lcd_i2c_cs_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_lcd_i2c_cs_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_lcd_i2c_cs_s1_end_xfer <= 1;
      else 
        d1_lcd_i2c_cs_s1_end_xfer <= lcd_i2c_cs_s1_end_xfer;
    end


  //lcd_i2c_cs_s1_waits_for_read in a cycle, which is an e_mux
  assign lcd_i2c_cs_s1_waits_for_read = lcd_i2c_cs_s1_in_a_read_cycle & lcd_i2c_cs_s1_begins_xfer;

  //lcd_i2c_cs_s1_in_a_read_cycle assignment, which is an e_assign
  assign lcd_i2c_cs_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = lcd_i2c_cs_s1_in_a_read_cycle;

  //lcd_i2c_cs_s1_waits_for_write in a cycle, which is an e_mux
  assign lcd_i2c_cs_s1_waits_for_write = lcd_i2c_cs_s1_in_a_write_cycle & 0;

  //lcd_i2c_cs_s1_in_a_write_cycle assignment, which is an e_assign
  assign lcd_i2c_cs_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = lcd_i2c_cs_s1_in_a_write_cycle;

  assign wait_for_lcd_i2c_cs_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_i2c_cs/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_i2c_dat_s1_arbitrator (
                                   // inputs:
                                    clk,
                                    clock_crossing_bridge_m1_address_to_slave,
                                    clock_crossing_bridge_m1_latency_counter,
                                    clock_crossing_bridge_m1_nativeaddress,
                                    clock_crossing_bridge_m1_read,
                                    clock_crossing_bridge_m1_write,
                                    clock_crossing_bridge_m1_writedata,
                                    lcd_i2c_dat_s1_readdata,
                                    reset_n,

                                   // outputs:
                                    clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1,
                                    clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1,
                                    clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1,
                                    clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1,
                                    d1_lcd_i2c_dat_s1_end_xfer,
                                    lcd_i2c_dat_s1_address,
                                    lcd_i2c_dat_s1_chipselect,
                                    lcd_i2c_dat_s1_readdata_from_sa,
                                    lcd_i2c_dat_s1_reset_n,
                                    lcd_i2c_dat_s1_write_n,
                                    lcd_i2c_dat_s1_writedata
                                 )
;

  output           clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1;
  output           clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1;
  output           clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1;
  output           clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1;
  output           d1_lcd_i2c_dat_s1_end_xfer;
  output  [  1: 0] lcd_i2c_dat_s1_address;
  output           lcd_i2c_dat_s1_chipselect;
  output  [ 31: 0] lcd_i2c_dat_s1_readdata_from_sa;
  output           lcd_i2c_dat_s1_reset_n;
  output           lcd_i2c_dat_s1_write_n;
  output  [ 31: 0] lcd_i2c_dat_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] lcd_i2c_dat_s1_readdata;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_saved_grant_lcd_i2c_dat_s1;
  reg              d1_lcd_i2c_dat_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_lcd_i2c_dat_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] lcd_i2c_dat_s1_address;
  wire             lcd_i2c_dat_s1_allgrants;
  wire             lcd_i2c_dat_s1_allow_new_arb_cycle;
  wire             lcd_i2c_dat_s1_any_bursting_master_saved_grant;
  wire             lcd_i2c_dat_s1_any_continuerequest;
  wire             lcd_i2c_dat_s1_arb_counter_enable;
  reg              lcd_i2c_dat_s1_arb_share_counter;
  wire             lcd_i2c_dat_s1_arb_share_counter_next_value;
  wire             lcd_i2c_dat_s1_arb_share_set_values;
  wire             lcd_i2c_dat_s1_beginbursttransfer_internal;
  wire             lcd_i2c_dat_s1_begins_xfer;
  wire             lcd_i2c_dat_s1_chipselect;
  wire             lcd_i2c_dat_s1_end_xfer;
  wire             lcd_i2c_dat_s1_firsttransfer;
  wire             lcd_i2c_dat_s1_grant_vector;
  wire             lcd_i2c_dat_s1_in_a_read_cycle;
  wire             lcd_i2c_dat_s1_in_a_write_cycle;
  wire             lcd_i2c_dat_s1_master_qreq_vector;
  wire             lcd_i2c_dat_s1_non_bursting_master_requests;
  wire    [ 31: 0] lcd_i2c_dat_s1_readdata_from_sa;
  reg              lcd_i2c_dat_s1_reg_firsttransfer;
  wire             lcd_i2c_dat_s1_reset_n;
  reg              lcd_i2c_dat_s1_slavearbiterlockenable;
  wire             lcd_i2c_dat_s1_slavearbiterlockenable2;
  wire             lcd_i2c_dat_s1_unreg_firsttransfer;
  wire             lcd_i2c_dat_s1_waits_for_read;
  wire             lcd_i2c_dat_s1_waits_for_write;
  wire             lcd_i2c_dat_s1_write_n;
  wire    [ 31: 0] lcd_i2c_dat_s1_writedata;
  wire             wait_for_lcd_i2c_dat_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~lcd_i2c_dat_s1_end_xfer;
    end


  assign lcd_i2c_dat_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1));
  //assign lcd_i2c_dat_s1_readdata_from_sa = lcd_i2c_dat_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_i2c_dat_s1_readdata_from_sa = lcd_i2c_dat_s1_readdata;

  assign clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h400) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //lcd_i2c_dat_s1_arb_share_counter set values, which is an e_mux
  assign lcd_i2c_dat_s1_arb_share_set_values = 1;

  //lcd_i2c_dat_s1_non_bursting_master_requests mux, which is an e_mux
  assign lcd_i2c_dat_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1;

  //lcd_i2c_dat_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign lcd_i2c_dat_s1_any_bursting_master_saved_grant = 0;

  //lcd_i2c_dat_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign lcd_i2c_dat_s1_arb_share_counter_next_value = lcd_i2c_dat_s1_firsttransfer ? (lcd_i2c_dat_s1_arb_share_set_values - 1) : |lcd_i2c_dat_s1_arb_share_counter ? (lcd_i2c_dat_s1_arb_share_counter - 1) : 0;

  //lcd_i2c_dat_s1_allgrants all slave grants, which is an e_mux
  assign lcd_i2c_dat_s1_allgrants = |lcd_i2c_dat_s1_grant_vector;

  //lcd_i2c_dat_s1_end_xfer assignment, which is an e_assign
  assign lcd_i2c_dat_s1_end_xfer = ~(lcd_i2c_dat_s1_waits_for_read | lcd_i2c_dat_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_lcd_i2c_dat_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_lcd_i2c_dat_s1 = lcd_i2c_dat_s1_end_xfer & (~lcd_i2c_dat_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //lcd_i2c_dat_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign lcd_i2c_dat_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_lcd_i2c_dat_s1 & lcd_i2c_dat_s1_allgrants) | (end_xfer_arb_share_counter_term_lcd_i2c_dat_s1 & ~lcd_i2c_dat_s1_non_bursting_master_requests);

  //lcd_i2c_dat_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_dat_s1_arb_share_counter <= 0;
      else if (lcd_i2c_dat_s1_arb_counter_enable)
          lcd_i2c_dat_s1_arb_share_counter <= lcd_i2c_dat_s1_arb_share_counter_next_value;
    end


  //lcd_i2c_dat_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_dat_s1_slavearbiterlockenable <= 0;
      else if ((|lcd_i2c_dat_s1_master_qreq_vector & end_xfer_arb_share_counter_term_lcd_i2c_dat_s1) | (end_xfer_arb_share_counter_term_lcd_i2c_dat_s1 & ~lcd_i2c_dat_s1_non_bursting_master_requests))
          lcd_i2c_dat_s1_slavearbiterlockenable <= |lcd_i2c_dat_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 lcd_i2c_dat/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = lcd_i2c_dat_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //lcd_i2c_dat_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign lcd_i2c_dat_s1_slavearbiterlockenable2 = |lcd_i2c_dat_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 lcd_i2c_dat/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = lcd_i2c_dat_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //lcd_i2c_dat_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign lcd_i2c_dat_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1 = clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1 = clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1 & clock_crossing_bridge_m1_read & ~lcd_i2c_dat_s1_waits_for_read;

  //lcd_i2c_dat_s1_writedata mux, which is an e_mux
  assign lcd_i2c_dat_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1 = clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1;

  //clock_crossing_bridge/m1 saved-grant lcd_i2c_dat/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_lcd_i2c_dat_s1 = clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1;

  //allow new arb cycle for lcd_i2c_dat/s1, which is an e_assign
  assign lcd_i2c_dat_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign lcd_i2c_dat_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign lcd_i2c_dat_s1_master_qreq_vector = 1;

  //lcd_i2c_dat_s1_reset_n assignment, which is an e_assign
  assign lcd_i2c_dat_s1_reset_n = reset_n;

  assign lcd_i2c_dat_s1_chipselect = clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1;
  //lcd_i2c_dat_s1_firsttransfer first transaction, which is an e_assign
  assign lcd_i2c_dat_s1_firsttransfer = lcd_i2c_dat_s1_begins_xfer ? lcd_i2c_dat_s1_unreg_firsttransfer : lcd_i2c_dat_s1_reg_firsttransfer;

  //lcd_i2c_dat_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign lcd_i2c_dat_s1_unreg_firsttransfer = ~(lcd_i2c_dat_s1_slavearbiterlockenable & lcd_i2c_dat_s1_any_continuerequest);

  //lcd_i2c_dat_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_dat_s1_reg_firsttransfer <= 1'b1;
      else if (lcd_i2c_dat_s1_begins_xfer)
          lcd_i2c_dat_s1_reg_firsttransfer <= lcd_i2c_dat_s1_unreg_firsttransfer;
    end


  //lcd_i2c_dat_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign lcd_i2c_dat_s1_beginbursttransfer_internal = lcd_i2c_dat_s1_begins_xfer;

  //~lcd_i2c_dat_s1_write_n assignment, which is an e_mux
  assign lcd_i2c_dat_s1_write_n = ~(clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1 & clock_crossing_bridge_m1_write);

  //lcd_i2c_dat_s1_address mux, which is an e_mux
  assign lcd_i2c_dat_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_lcd_i2c_dat_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_lcd_i2c_dat_s1_end_xfer <= 1;
      else 
        d1_lcd_i2c_dat_s1_end_xfer <= lcd_i2c_dat_s1_end_xfer;
    end


  //lcd_i2c_dat_s1_waits_for_read in a cycle, which is an e_mux
  assign lcd_i2c_dat_s1_waits_for_read = lcd_i2c_dat_s1_in_a_read_cycle & lcd_i2c_dat_s1_begins_xfer;

  //lcd_i2c_dat_s1_in_a_read_cycle assignment, which is an e_assign
  assign lcd_i2c_dat_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = lcd_i2c_dat_s1_in_a_read_cycle;

  //lcd_i2c_dat_s1_waits_for_write in a cycle, which is an e_mux
  assign lcd_i2c_dat_s1_waits_for_write = lcd_i2c_dat_s1_in_a_write_cycle & 0;

  //lcd_i2c_dat_s1_in_a_write_cycle assignment, which is an e_assign
  assign lcd_i2c_dat_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = lcd_i2c_dat_s1_in_a_write_cycle;

  assign wait_for_lcd_i2c_dat_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_i2c_dat/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_i2c_scl_s1_arbitrator (
                                   // inputs:
                                    clk,
                                    clock_crossing_bridge_m1_address_to_slave,
                                    clock_crossing_bridge_m1_latency_counter,
                                    clock_crossing_bridge_m1_nativeaddress,
                                    clock_crossing_bridge_m1_read,
                                    clock_crossing_bridge_m1_write,
                                    clock_crossing_bridge_m1_writedata,
                                    lcd_i2c_scl_s1_readdata,
                                    reset_n,

                                   // outputs:
                                    clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1,
                                    clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1,
                                    clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1,
                                    clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1,
                                    d1_lcd_i2c_scl_s1_end_xfer,
                                    lcd_i2c_scl_s1_address,
                                    lcd_i2c_scl_s1_chipselect,
                                    lcd_i2c_scl_s1_readdata_from_sa,
                                    lcd_i2c_scl_s1_reset_n,
                                    lcd_i2c_scl_s1_write_n,
                                    lcd_i2c_scl_s1_writedata
                                 )
;

  output           clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1;
  output           clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1;
  output           clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1;
  output           clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1;
  output           d1_lcd_i2c_scl_s1_end_xfer;
  output  [  1: 0] lcd_i2c_scl_s1_address;
  output           lcd_i2c_scl_s1_chipselect;
  output  [ 31: 0] lcd_i2c_scl_s1_readdata_from_sa;
  output           lcd_i2c_scl_s1_reset_n;
  output           lcd_i2c_scl_s1_write_n;
  output  [ 31: 0] lcd_i2c_scl_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] lcd_i2c_scl_s1_readdata;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_saved_grant_lcd_i2c_scl_s1;
  reg              d1_lcd_i2c_scl_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_lcd_i2c_scl_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] lcd_i2c_scl_s1_address;
  wire             lcd_i2c_scl_s1_allgrants;
  wire             lcd_i2c_scl_s1_allow_new_arb_cycle;
  wire             lcd_i2c_scl_s1_any_bursting_master_saved_grant;
  wire             lcd_i2c_scl_s1_any_continuerequest;
  wire             lcd_i2c_scl_s1_arb_counter_enable;
  reg              lcd_i2c_scl_s1_arb_share_counter;
  wire             lcd_i2c_scl_s1_arb_share_counter_next_value;
  wire             lcd_i2c_scl_s1_arb_share_set_values;
  wire             lcd_i2c_scl_s1_beginbursttransfer_internal;
  wire             lcd_i2c_scl_s1_begins_xfer;
  wire             lcd_i2c_scl_s1_chipselect;
  wire             lcd_i2c_scl_s1_end_xfer;
  wire             lcd_i2c_scl_s1_firsttransfer;
  wire             lcd_i2c_scl_s1_grant_vector;
  wire             lcd_i2c_scl_s1_in_a_read_cycle;
  wire             lcd_i2c_scl_s1_in_a_write_cycle;
  wire             lcd_i2c_scl_s1_master_qreq_vector;
  wire             lcd_i2c_scl_s1_non_bursting_master_requests;
  wire    [ 31: 0] lcd_i2c_scl_s1_readdata_from_sa;
  reg              lcd_i2c_scl_s1_reg_firsttransfer;
  wire             lcd_i2c_scl_s1_reset_n;
  reg              lcd_i2c_scl_s1_slavearbiterlockenable;
  wire             lcd_i2c_scl_s1_slavearbiterlockenable2;
  wire             lcd_i2c_scl_s1_unreg_firsttransfer;
  wire             lcd_i2c_scl_s1_waits_for_read;
  wire             lcd_i2c_scl_s1_waits_for_write;
  wire             lcd_i2c_scl_s1_write_n;
  wire    [ 31: 0] lcd_i2c_scl_s1_writedata;
  wire             wait_for_lcd_i2c_scl_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~lcd_i2c_scl_s1_end_xfer;
    end


  assign lcd_i2c_scl_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1));
  //assign lcd_i2c_scl_s1_readdata_from_sa = lcd_i2c_scl_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_i2c_scl_s1_readdata_from_sa = lcd_i2c_scl_s1_readdata;

  assign clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h300) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //lcd_i2c_scl_s1_arb_share_counter set values, which is an e_mux
  assign lcd_i2c_scl_s1_arb_share_set_values = 1;

  //lcd_i2c_scl_s1_non_bursting_master_requests mux, which is an e_mux
  assign lcd_i2c_scl_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1;

  //lcd_i2c_scl_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign lcd_i2c_scl_s1_any_bursting_master_saved_grant = 0;

  //lcd_i2c_scl_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign lcd_i2c_scl_s1_arb_share_counter_next_value = lcd_i2c_scl_s1_firsttransfer ? (lcd_i2c_scl_s1_arb_share_set_values - 1) : |lcd_i2c_scl_s1_arb_share_counter ? (lcd_i2c_scl_s1_arb_share_counter - 1) : 0;

  //lcd_i2c_scl_s1_allgrants all slave grants, which is an e_mux
  assign lcd_i2c_scl_s1_allgrants = |lcd_i2c_scl_s1_grant_vector;

  //lcd_i2c_scl_s1_end_xfer assignment, which is an e_assign
  assign lcd_i2c_scl_s1_end_xfer = ~(lcd_i2c_scl_s1_waits_for_read | lcd_i2c_scl_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 = lcd_i2c_scl_s1_end_xfer & (~lcd_i2c_scl_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //lcd_i2c_scl_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign lcd_i2c_scl_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 & lcd_i2c_scl_s1_allgrants) | (end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 & ~lcd_i2c_scl_s1_non_bursting_master_requests);

  //lcd_i2c_scl_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_scl_s1_arb_share_counter <= 0;
      else if (lcd_i2c_scl_s1_arb_counter_enable)
          lcd_i2c_scl_s1_arb_share_counter <= lcd_i2c_scl_s1_arb_share_counter_next_value;
    end


  //lcd_i2c_scl_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_scl_s1_slavearbiterlockenable <= 0;
      else if ((|lcd_i2c_scl_s1_master_qreq_vector & end_xfer_arb_share_counter_term_lcd_i2c_scl_s1) | (end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 & ~lcd_i2c_scl_s1_non_bursting_master_requests))
          lcd_i2c_scl_s1_slavearbiterlockenable <= |lcd_i2c_scl_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 lcd_i2c_scl/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = lcd_i2c_scl_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //lcd_i2c_scl_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign lcd_i2c_scl_s1_slavearbiterlockenable2 = |lcd_i2c_scl_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 lcd_i2c_scl/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = lcd_i2c_scl_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //lcd_i2c_scl_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign lcd_i2c_scl_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1 = clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1 = clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1 & clock_crossing_bridge_m1_read & ~lcd_i2c_scl_s1_waits_for_read;

  //lcd_i2c_scl_s1_writedata mux, which is an e_mux
  assign lcd_i2c_scl_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1 = clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1;

  //clock_crossing_bridge/m1 saved-grant lcd_i2c_scl/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_lcd_i2c_scl_s1 = clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1;

  //allow new arb cycle for lcd_i2c_scl/s1, which is an e_assign
  assign lcd_i2c_scl_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign lcd_i2c_scl_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign lcd_i2c_scl_s1_master_qreq_vector = 1;

  //lcd_i2c_scl_s1_reset_n assignment, which is an e_assign
  assign lcd_i2c_scl_s1_reset_n = reset_n;

  assign lcd_i2c_scl_s1_chipselect = clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1;
  //lcd_i2c_scl_s1_firsttransfer first transaction, which is an e_assign
  assign lcd_i2c_scl_s1_firsttransfer = lcd_i2c_scl_s1_begins_xfer ? lcd_i2c_scl_s1_unreg_firsttransfer : lcd_i2c_scl_s1_reg_firsttransfer;

  //lcd_i2c_scl_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign lcd_i2c_scl_s1_unreg_firsttransfer = ~(lcd_i2c_scl_s1_slavearbiterlockenable & lcd_i2c_scl_s1_any_continuerequest);

  //lcd_i2c_scl_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_i2c_scl_s1_reg_firsttransfer <= 1'b1;
      else if (lcd_i2c_scl_s1_begins_xfer)
          lcd_i2c_scl_s1_reg_firsttransfer <= lcd_i2c_scl_s1_unreg_firsttransfer;
    end


  //lcd_i2c_scl_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign lcd_i2c_scl_s1_beginbursttransfer_internal = lcd_i2c_scl_s1_begins_xfer;

  //~lcd_i2c_scl_s1_write_n assignment, which is an e_mux
  assign lcd_i2c_scl_s1_write_n = ~(clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1 & clock_crossing_bridge_m1_write);

  //lcd_i2c_scl_s1_address mux, which is an e_mux
  assign lcd_i2c_scl_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_lcd_i2c_scl_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_lcd_i2c_scl_s1_end_xfer <= 1;
      else 
        d1_lcd_i2c_scl_s1_end_xfer <= lcd_i2c_scl_s1_end_xfer;
    end


  //lcd_i2c_scl_s1_waits_for_read in a cycle, which is an e_mux
  assign lcd_i2c_scl_s1_waits_for_read = lcd_i2c_scl_s1_in_a_read_cycle & lcd_i2c_scl_s1_begins_xfer;

  //lcd_i2c_scl_s1_in_a_read_cycle assignment, which is an e_assign
  assign lcd_i2c_scl_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = lcd_i2c_scl_s1_in_a_read_cycle;

  //lcd_i2c_scl_s1_waits_for_write in a cycle, which is an e_mux
  assign lcd_i2c_scl_s1_waits_for_write = lcd_i2c_scl_s1_in_a_write_cycle & 0;

  //lcd_i2c_scl_s1_in_a_write_cycle assignment, which is an e_assign
  assign lcd_i2c_scl_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = lcd_i2c_scl_s1_in_a_write_cycle;

  assign wait_for_lcd_i2c_scl_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_i2c_scl/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_on_chip_memory_fifo_in_arbitrator (
                                               // inputs:
                                                clk,
                                                lcd_on_chip_memory_fifo_in_ready,
                                                lcd_ta_formatter_to_fifo_out_data,
                                                lcd_ta_formatter_to_fifo_out_endofpacket,
                                                lcd_ta_formatter_to_fifo_out_startofpacket,
                                                lcd_ta_formatter_to_fifo_out_valid,
                                                reset_n,

                                               // outputs:
                                                lcd_on_chip_memory_fifo_in_data,
                                                lcd_on_chip_memory_fifo_in_endofpacket,
                                                lcd_on_chip_memory_fifo_in_ready_from_sa,
                                                lcd_on_chip_memory_fifo_in_reset_n,
                                                lcd_on_chip_memory_fifo_in_startofpacket,
                                                lcd_on_chip_memory_fifo_in_valid
                                             )
;

  output  [  7: 0] lcd_on_chip_memory_fifo_in_data;
  output           lcd_on_chip_memory_fifo_in_endofpacket;
  output           lcd_on_chip_memory_fifo_in_ready_from_sa;
  output           lcd_on_chip_memory_fifo_in_reset_n;
  output           lcd_on_chip_memory_fifo_in_startofpacket;
  output           lcd_on_chip_memory_fifo_in_valid;
  input            clk;
  input            lcd_on_chip_memory_fifo_in_ready;
  input   [  7: 0] lcd_ta_formatter_to_fifo_out_data;
  input            lcd_ta_formatter_to_fifo_out_endofpacket;
  input            lcd_ta_formatter_to_fifo_out_startofpacket;
  input            lcd_ta_formatter_to_fifo_out_valid;
  input            reset_n;

  wire    [  7: 0] lcd_on_chip_memory_fifo_in_data;
  wire             lcd_on_chip_memory_fifo_in_endofpacket;
  wire             lcd_on_chip_memory_fifo_in_ready_from_sa;
  wire             lcd_on_chip_memory_fifo_in_reset_n;
  wire             lcd_on_chip_memory_fifo_in_startofpacket;
  wire             lcd_on_chip_memory_fifo_in_valid;
  //mux lcd_on_chip_memory_fifo_in_data, which is an e_mux
  assign lcd_on_chip_memory_fifo_in_data = lcd_ta_formatter_to_fifo_out_data;

  //mux lcd_on_chip_memory_fifo_in_endofpacket, which is an e_mux
  assign lcd_on_chip_memory_fifo_in_endofpacket = lcd_ta_formatter_to_fifo_out_endofpacket;

  //assign lcd_on_chip_memory_fifo_in_ready_from_sa = lcd_on_chip_memory_fifo_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_on_chip_memory_fifo_in_ready_from_sa = lcd_on_chip_memory_fifo_in_ready;

  //mux lcd_on_chip_memory_fifo_in_startofpacket, which is an e_mux
  assign lcd_on_chip_memory_fifo_in_startofpacket = lcd_ta_formatter_to_fifo_out_startofpacket;

  //mux lcd_on_chip_memory_fifo_in_valid, which is an e_mux
  assign lcd_on_chip_memory_fifo_in_valid = lcd_ta_formatter_to_fifo_out_valid;

  //lcd_on_chip_memory_fifo_in_reset_n assignment, which is an e_assign
  assign lcd_on_chip_memory_fifo_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_on_chip_memory_fifo_out_arbitrator (
                                                // inputs:
                                                 clk,
                                                 lcd_on_chip_memory_fifo_out_data,
                                                 lcd_on_chip_memory_fifo_out_endofpacket,
                                                 lcd_on_chip_memory_fifo_out_startofpacket,
                                                 lcd_on_chip_memory_fifo_out_valid,
                                                 lcd_ta_fifo_to_sequencer_in_ready_from_sa,
                                                 reset_n,

                                                // outputs:
                                                 lcd_on_chip_memory_fifo_out_ready,
                                                 lcd_on_chip_memory_fifo_out_reset_n
                                              )
;

  output           lcd_on_chip_memory_fifo_out_ready;
  output           lcd_on_chip_memory_fifo_out_reset_n;
  input            clk;
  input   [  7: 0] lcd_on_chip_memory_fifo_out_data;
  input            lcd_on_chip_memory_fifo_out_endofpacket;
  input            lcd_on_chip_memory_fifo_out_startofpacket;
  input            lcd_on_chip_memory_fifo_out_valid;
  input            lcd_ta_fifo_to_sequencer_in_ready_from_sa;
  input            reset_n;

  wire             lcd_on_chip_memory_fifo_out_ready;
  wire             lcd_on_chip_memory_fifo_out_reset_n;
  //lcd_on_chip_memory_fifo_out_reset_n assignment, which is an e_assign
  assign lcd_on_chip_memory_fifo_out_reset_n = reset_n;

  //mux lcd_on_chip_memory_fifo_out_ready, which is an e_mux
  assign lcd_on_chip_memory_fifo_out_ready = lcd_ta_fifo_to_sequencer_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_pixel_converter_in_arbitrator (
                                           // inputs:
                                            clk,
                                            lcd_pixel_converter_in_ready,
                                            lcd_sgdma_out_data,
                                            lcd_sgdma_out_empty,
                                            lcd_sgdma_out_endofpacket,
                                            lcd_sgdma_out_startofpacket,
                                            lcd_sgdma_out_valid,
                                            reset_n,

                                           // outputs:
                                            lcd_pixel_converter_in_data,
                                            lcd_pixel_converter_in_empty,
                                            lcd_pixel_converter_in_endofpacket,
                                            lcd_pixel_converter_in_ready_from_sa,
                                            lcd_pixel_converter_in_reset_n,
                                            lcd_pixel_converter_in_startofpacket,
                                            lcd_pixel_converter_in_valid
                                         )
;

  output  [ 31: 0] lcd_pixel_converter_in_data;
  output  [  1: 0] lcd_pixel_converter_in_empty;
  output           lcd_pixel_converter_in_endofpacket;
  output           lcd_pixel_converter_in_ready_from_sa;
  output           lcd_pixel_converter_in_reset_n;
  output           lcd_pixel_converter_in_startofpacket;
  output           lcd_pixel_converter_in_valid;
  input            clk;
  input            lcd_pixel_converter_in_ready;
  input   [ 31: 0] lcd_sgdma_out_data;
  input   [  1: 0] lcd_sgdma_out_empty;
  input            lcd_sgdma_out_endofpacket;
  input            lcd_sgdma_out_startofpacket;
  input            lcd_sgdma_out_valid;
  input            reset_n;

  wire    [ 31: 0] lcd_pixel_converter_in_data;
  wire    [  1: 0] lcd_pixel_converter_in_empty;
  wire             lcd_pixel_converter_in_endofpacket;
  wire             lcd_pixel_converter_in_ready_from_sa;
  wire             lcd_pixel_converter_in_reset_n;
  wire             lcd_pixel_converter_in_startofpacket;
  wire             lcd_pixel_converter_in_valid;
  //mux lcd_pixel_converter_in_data, which is an e_mux
  assign lcd_pixel_converter_in_data = lcd_sgdma_out_data;

  //mux lcd_pixel_converter_in_empty, which is an e_mux
  assign lcd_pixel_converter_in_empty = lcd_sgdma_out_empty;

  //mux lcd_pixel_converter_in_endofpacket, which is an e_mux
  assign lcd_pixel_converter_in_endofpacket = lcd_sgdma_out_endofpacket;

  //assign lcd_pixel_converter_in_ready_from_sa = lcd_pixel_converter_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_pixel_converter_in_ready_from_sa = lcd_pixel_converter_in_ready;

  //mux lcd_pixel_converter_in_startofpacket, which is an e_mux
  assign lcd_pixel_converter_in_startofpacket = lcd_sgdma_out_startofpacket;

  //mux lcd_pixel_converter_in_valid, which is an e_mux
  assign lcd_pixel_converter_in_valid = lcd_sgdma_out_valid;

  //lcd_pixel_converter_in_reset_n assignment, which is an e_assign
  assign lcd_pixel_converter_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_pixel_converter_out_arbitrator (
                                            // inputs:
                                             clk,
                                             lcd_data_format_adapter_in_ready_from_sa,
                                             lcd_pixel_converter_out_data,
                                             lcd_pixel_converter_out_empty,
                                             lcd_pixel_converter_out_endofpacket,
                                             lcd_pixel_converter_out_startofpacket,
                                             lcd_pixel_converter_out_valid,
                                             reset_n,

                                            // outputs:
                                             lcd_pixel_converter_out_ready
                                          )
;

  output           lcd_pixel_converter_out_ready;
  input            clk;
  input            lcd_data_format_adapter_in_ready_from_sa;
  input   [ 23: 0] lcd_pixel_converter_out_data;
  input   [  1: 0] lcd_pixel_converter_out_empty;
  input            lcd_pixel_converter_out_endofpacket;
  input            lcd_pixel_converter_out_startofpacket;
  input            lcd_pixel_converter_out_valid;
  input            reset_n;

  wire             lcd_pixel_converter_out_ready;
  //mux lcd_pixel_converter_out_ready, which is an e_mux
  assign lcd_pixel_converter_out_ready = lcd_data_format_adapter_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_sgdma_csr_arbitrator (
                                  // inputs:
                                   clk,
                                   lcd_sgdma_csr_irq,
                                   lcd_sgdma_csr_readdata,
                                   pipeline_bridge_m1_address_to_slave,
                                   pipeline_bridge_m1_burstcount,
                                   pipeline_bridge_m1_chipselect,
                                   pipeline_bridge_m1_latency_counter,
                                   pipeline_bridge_m1_read,
                                   pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                   pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                   pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                   pipeline_bridge_m1_write,
                                   pipeline_bridge_m1_writedata,
                                   reset_n,

                                  // outputs:
                                   d1_lcd_sgdma_csr_end_xfer,
                                   lcd_sgdma_csr_address,
                                   lcd_sgdma_csr_chipselect,
                                   lcd_sgdma_csr_irq_from_sa,
                                   lcd_sgdma_csr_read,
                                   lcd_sgdma_csr_readdata_from_sa,
                                   lcd_sgdma_csr_reset_n,
                                   lcd_sgdma_csr_write,
                                   lcd_sgdma_csr_writedata,
                                   pipeline_bridge_m1_granted_lcd_sgdma_csr,
                                   pipeline_bridge_m1_qualified_request_lcd_sgdma_csr,
                                   pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr,
                                   pipeline_bridge_m1_requests_lcd_sgdma_csr
                                )
;

  output           d1_lcd_sgdma_csr_end_xfer;
  output  [  3: 0] lcd_sgdma_csr_address;
  output           lcd_sgdma_csr_chipselect;
  output           lcd_sgdma_csr_irq_from_sa;
  output           lcd_sgdma_csr_read;
  output  [ 31: 0] lcd_sgdma_csr_readdata_from_sa;
  output           lcd_sgdma_csr_reset_n;
  output           lcd_sgdma_csr_write;
  output  [ 31: 0] lcd_sgdma_csr_writedata;
  output           pipeline_bridge_m1_granted_lcd_sgdma_csr;
  output           pipeline_bridge_m1_qualified_request_lcd_sgdma_csr;
  output           pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr;
  output           pipeline_bridge_m1_requests_lcd_sgdma_csr;
  input            clk;
  input            lcd_sgdma_csr_irq;
  input   [ 31: 0] lcd_sgdma_csr_readdata;
  input   [ 26: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              d1_lcd_sgdma_csr_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_lcd_sgdma_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  3: 0] lcd_sgdma_csr_address;
  wire             lcd_sgdma_csr_allgrants;
  wire             lcd_sgdma_csr_allow_new_arb_cycle;
  wire             lcd_sgdma_csr_any_bursting_master_saved_grant;
  wire             lcd_sgdma_csr_any_continuerequest;
  wire             lcd_sgdma_csr_arb_counter_enable;
  reg              lcd_sgdma_csr_arb_share_counter;
  wire             lcd_sgdma_csr_arb_share_counter_next_value;
  wire             lcd_sgdma_csr_arb_share_set_values;
  wire             lcd_sgdma_csr_beginbursttransfer_internal;
  wire             lcd_sgdma_csr_begins_xfer;
  wire             lcd_sgdma_csr_chipselect;
  wire             lcd_sgdma_csr_end_xfer;
  wire             lcd_sgdma_csr_firsttransfer;
  wire             lcd_sgdma_csr_grant_vector;
  wire             lcd_sgdma_csr_in_a_read_cycle;
  wire             lcd_sgdma_csr_in_a_write_cycle;
  wire             lcd_sgdma_csr_irq_from_sa;
  wire             lcd_sgdma_csr_master_qreq_vector;
  wire             lcd_sgdma_csr_non_bursting_master_requests;
  wire             lcd_sgdma_csr_read;
  wire    [ 31: 0] lcd_sgdma_csr_readdata_from_sa;
  reg              lcd_sgdma_csr_reg_firsttransfer;
  wire             lcd_sgdma_csr_reset_n;
  reg              lcd_sgdma_csr_slavearbiterlockenable;
  wire             lcd_sgdma_csr_slavearbiterlockenable2;
  wire             lcd_sgdma_csr_unreg_firsttransfer;
  wire             lcd_sgdma_csr_waits_for_read;
  wire             lcd_sgdma_csr_waits_for_write;
  wire             lcd_sgdma_csr_write;
  wire    [ 31: 0] lcd_sgdma_csr_writedata;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_qualified_request_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_requests_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_saved_grant_lcd_sgdma_csr;
  wire    [ 26: 0] shifted_address_to_lcd_sgdma_csr_from_pipeline_bridge_m1;
  wire             wait_for_lcd_sgdma_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~lcd_sgdma_csr_end_xfer;
    end


  assign lcd_sgdma_csr_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_lcd_sgdma_csr));
  //assign lcd_sgdma_csr_readdata_from_sa = lcd_sgdma_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_sgdma_csr_readdata_from_sa = lcd_sgdma_csr_readdata;

  assign pipeline_bridge_m1_requests_lcd_sgdma_csr = ({pipeline_bridge_m1_address_to_slave[26 : 6] , 6'b0} == 27'h4401800) & pipeline_bridge_m1_chipselect;
  //lcd_sgdma_csr_arb_share_counter set values, which is an e_mux
  assign lcd_sgdma_csr_arb_share_set_values = 1;

  //lcd_sgdma_csr_non_bursting_master_requests mux, which is an e_mux
  assign lcd_sgdma_csr_non_bursting_master_requests = pipeline_bridge_m1_requests_lcd_sgdma_csr;

  //lcd_sgdma_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign lcd_sgdma_csr_any_bursting_master_saved_grant = 0;

  //lcd_sgdma_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign lcd_sgdma_csr_arb_share_counter_next_value = lcd_sgdma_csr_firsttransfer ? (lcd_sgdma_csr_arb_share_set_values - 1) : |lcd_sgdma_csr_arb_share_counter ? (lcd_sgdma_csr_arb_share_counter - 1) : 0;

  //lcd_sgdma_csr_allgrants all slave grants, which is an e_mux
  assign lcd_sgdma_csr_allgrants = |lcd_sgdma_csr_grant_vector;

  //lcd_sgdma_csr_end_xfer assignment, which is an e_assign
  assign lcd_sgdma_csr_end_xfer = ~(lcd_sgdma_csr_waits_for_read | lcd_sgdma_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_lcd_sgdma_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_lcd_sgdma_csr = lcd_sgdma_csr_end_xfer & (~lcd_sgdma_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //lcd_sgdma_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign lcd_sgdma_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_lcd_sgdma_csr & lcd_sgdma_csr_allgrants) | (end_xfer_arb_share_counter_term_lcd_sgdma_csr & ~lcd_sgdma_csr_non_bursting_master_requests);

  //lcd_sgdma_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_csr_arb_share_counter <= 0;
      else if (lcd_sgdma_csr_arb_counter_enable)
          lcd_sgdma_csr_arb_share_counter <= lcd_sgdma_csr_arb_share_counter_next_value;
    end


  //lcd_sgdma_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_csr_slavearbiterlockenable <= 0;
      else if ((|lcd_sgdma_csr_master_qreq_vector & end_xfer_arb_share_counter_term_lcd_sgdma_csr) | (end_xfer_arb_share_counter_term_lcd_sgdma_csr & ~lcd_sgdma_csr_non_bursting_master_requests))
          lcd_sgdma_csr_slavearbiterlockenable <= |lcd_sgdma_csr_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 lcd_sgdma/csr arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = lcd_sgdma_csr_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //lcd_sgdma_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign lcd_sgdma_csr_slavearbiterlockenable2 = |lcd_sgdma_csr_arb_share_counter_next_value;

  //pipeline_bridge/m1 lcd_sgdma/csr arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = lcd_sgdma_csr_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //lcd_sgdma_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign lcd_sgdma_csr_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_lcd_sgdma_csr = pipeline_bridge_m1_requests_lcd_sgdma_csr & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0) | (|pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register) | (|pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr = pipeline_bridge_m1_granted_lcd_sgdma_csr & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~lcd_sgdma_csr_waits_for_read;

  //lcd_sgdma_csr_writedata mux, which is an e_mux
  assign lcd_sgdma_csr_writedata = pipeline_bridge_m1_writedata;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_lcd_sgdma_csr = pipeline_bridge_m1_qualified_request_lcd_sgdma_csr;

  //pipeline_bridge/m1 saved-grant lcd_sgdma/csr, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_lcd_sgdma_csr = pipeline_bridge_m1_requests_lcd_sgdma_csr;

  //allow new arb cycle for lcd_sgdma/csr, which is an e_assign
  assign lcd_sgdma_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign lcd_sgdma_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign lcd_sgdma_csr_master_qreq_vector = 1;

  //lcd_sgdma_csr_reset_n assignment, which is an e_assign
  assign lcd_sgdma_csr_reset_n = reset_n;

  assign lcd_sgdma_csr_chipselect = pipeline_bridge_m1_granted_lcd_sgdma_csr;
  //lcd_sgdma_csr_firsttransfer first transaction, which is an e_assign
  assign lcd_sgdma_csr_firsttransfer = lcd_sgdma_csr_begins_xfer ? lcd_sgdma_csr_unreg_firsttransfer : lcd_sgdma_csr_reg_firsttransfer;

  //lcd_sgdma_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign lcd_sgdma_csr_unreg_firsttransfer = ~(lcd_sgdma_csr_slavearbiterlockenable & lcd_sgdma_csr_any_continuerequest);

  //lcd_sgdma_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_csr_reg_firsttransfer <= 1'b1;
      else if (lcd_sgdma_csr_begins_xfer)
          lcd_sgdma_csr_reg_firsttransfer <= lcd_sgdma_csr_unreg_firsttransfer;
    end


  //lcd_sgdma_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign lcd_sgdma_csr_beginbursttransfer_internal = lcd_sgdma_csr_begins_xfer;

  //lcd_sgdma_csr_read assignment, which is an e_mux
  assign lcd_sgdma_csr_read = pipeline_bridge_m1_granted_lcd_sgdma_csr & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //lcd_sgdma_csr_write assignment, which is an e_mux
  assign lcd_sgdma_csr_write = pipeline_bridge_m1_granted_lcd_sgdma_csr & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_lcd_sgdma_csr_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //lcd_sgdma_csr_address mux, which is an e_mux
  assign lcd_sgdma_csr_address = shifted_address_to_lcd_sgdma_csr_from_pipeline_bridge_m1 >> 2;

  //d1_lcd_sgdma_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_lcd_sgdma_csr_end_xfer <= 1;
      else 
        d1_lcd_sgdma_csr_end_xfer <= lcd_sgdma_csr_end_xfer;
    end


  //lcd_sgdma_csr_waits_for_read in a cycle, which is an e_mux
  assign lcd_sgdma_csr_waits_for_read = lcd_sgdma_csr_in_a_read_cycle & lcd_sgdma_csr_begins_xfer;

  //lcd_sgdma_csr_in_a_read_cycle assignment, which is an e_assign
  assign lcd_sgdma_csr_in_a_read_cycle = pipeline_bridge_m1_granted_lcd_sgdma_csr & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = lcd_sgdma_csr_in_a_read_cycle;

  //lcd_sgdma_csr_waits_for_write in a cycle, which is an e_mux
  assign lcd_sgdma_csr_waits_for_write = lcd_sgdma_csr_in_a_write_cycle & 0;

  //lcd_sgdma_csr_in_a_write_cycle assignment, which is an e_assign
  assign lcd_sgdma_csr_in_a_write_cycle = pipeline_bridge_m1_granted_lcd_sgdma_csr & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = lcd_sgdma_csr_in_a_write_cycle;

  assign wait_for_lcd_sgdma_csr_counter = 0;
  //assign lcd_sgdma_csr_irq_from_sa = lcd_sgdma_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_sgdma_csr_irq_from_sa = lcd_sgdma_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_sgdma/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_lcd_sgdma_csr && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave lcd_sgdma/csr", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_sgdma_descriptor_read_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_descriptor_memory_s2_end_xfer,
                                               descriptor_memory_s2_readdata_from_sa,
                                               lcd_sgdma_descriptor_read_address,
                                               lcd_sgdma_descriptor_read_granted_descriptor_memory_s2,
                                               lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2,
                                               lcd_sgdma_descriptor_read_read,
                                               lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2,
                                               lcd_sgdma_descriptor_read_requests_descriptor_memory_s2,
                                               reset_n,

                                              // outputs:
                                               lcd_sgdma_descriptor_read_address_to_slave,
                                               lcd_sgdma_descriptor_read_latency_counter,
                                               lcd_sgdma_descriptor_read_readdata,
                                               lcd_sgdma_descriptor_read_readdatavalid,
                                               lcd_sgdma_descriptor_read_waitrequest
                                            )
;

  output  [ 31: 0] lcd_sgdma_descriptor_read_address_to_slave;
  output           lcd_sgdma_descriptor_read_latency_counter;
  output  [ 31: 0] lcd_sgdma_descriptor_read_readdata;
  output           lcd_sgdma_descriptor_read_readdatavalid;
  output           lcd_sgdma_descriptor_read_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s2_end_xfer;
  input   [ 31: 0] descriptor_memory_s2_readdata_from_sa;
  input   [ 31: 0] lcd_sgdma_descriptor_read_address;
  input            lcd_sgdma_descriptor_read_granted_descriptor_memory_s2;
  input            lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2;
  input            lcd_sgdma_descriptor_read_read;
  input            lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2;
  input            lcd_sgdma_descriptor_read_requests_descriptor_memory_s2;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  reg     [ 31: 0] lcd_sgdma_descriptor_read_address_last_time;
  wire    [ 31: 0] lcd_sgdma_descriptor_read_address_to_slave;
  wire             lcd_sgdma_descriptor_read_is_granted_some_slave;
  reg              lcd_sgdma_descriptor_read_latency_counter;
  reg              lcd_sgdma_descriptor_read_read_but_no_slave_selected;
  reg              lcd_sgdma_descriptor_read_read_last_time;
  wire    [ 31: 0] lcd_sgdma_descriptor_read_readdata;
  wire             lcd_sgdma_descriptor_read_readdatavalid;
  wire             lcd_sgdma_descriptor_read_run;
  wire             lcd_sgdma_descriptor_read_waitrequest;
  wire             p1_lcd_sgdma_descriptor_read_latency_counter;
  wire             pre_flush_lcd_sgdma_descriptor_read_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2 | ~lcd_sgdma_descriptor_read_requests_descriptor_memory_s2) & (lcd_sgdma_descriptor_read_granted_descriptor_memory_s2 | ~lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2) & ((~lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2 | ~(lcd_sgdma_descriptor_read_read) | (1 & (lcd_sgdma_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign lcd_sgdma_descriptor_read_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign lcd_sgdma_descriptor_read_address_to_slave = {20'b100010000000000,
    lcd_sgdma_descriptor_read_address[11 : 0]};

  //lcd_sgdma_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        lcd_sgdma_descriptor_read_read_but_no_slave_selected <= lcd_sgdma_descriptor_read_read & lcd_sgdma_descriptor_read_run & ~lcd_sgdma_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign lcd_sgdma_descriptor_read_is_granted_some_slave = lcd_sgdma_descriptor_read_granted_descriptor_memory_s2;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_lcd_sgdma_descriptor_read_readdatavalid = lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign lcd_sgdma_descriptor_read_readdatavalid = lcd_sgdma_descriptor_read_read_but_no_slave_selected |
    pre_flush_lcd_sgdma_descriptor_read_readdatavalid;

  //lcd_sgdma/descriptor_read readdata mux, which is an e_mux
  assign lcd_sgdma_descriptor_read_readdata = descriptor_memory_s2_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign lcd_sgdma_descriptor_read_waitrequest = ~lcd_sgdma_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_read_latency_counter <= 0;
      else 
        lcd_sgdma_descriptor_read_latency_counter <= p1_lcd_sgdma_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_lcd_sgdma_descriptor_read_latency_counter = ((lcd_sgdma_descriptor_read_run & lcd_sgdma_descriptor_read_read))? latency_load_value :
    (lcd_sgdma_descriptor_read_latency_counter)? lcd_sgdma_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {lcd_sgdma_descriptor_read_requests_descriptor_memory_s2}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_sgdma_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_read_address_last_time <= 0;
      else 
        lcd_sgdma_descriptor_read_address_last_time <= lcd_sgdma_descriptor_read_address;
    end


  //lcd_sgdma/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= lcd_sgdma_descriptor_read_waitrequest & (lcd_sgdma_descriptor_read_read);
    end


  //lcd_sgdma_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_descriptor_read_address != lcd_sgdma_descriptor_read_address_last_time))
        begin
          $write("%0d ns: lcd_sgdma_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //lcd_sgdma_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_read_read_last_time <= 0;
      else 
        lcd_sgdma_descriptor_read_read_last_time <= lcd_sgdma_descriptor_read_read;
    end


  //lcd_sgdma_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_descriptor_read_read != lcd_sgdma_descriptor_read_read_last_time))
        begin
          $write("%0d ns: lcd_sgdma_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_sgdma_descriptor_write_arbitrator (
                                               // inputs:
                                                clk,
                                                d1_descriptor_memory_s2_end_xfer,
                                                lcd_sgdma_descriptor_write_address,
                                                lcd_sgdma_descriptor_write_granted_descriptor_memory_s2,
                                                lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2,
                                                lcd_sgdma_descriptor_write_requests_descriptor_memory_s2,
                                                lcd_sgdma_descriptor_write_write,
                                                lcd_sgdma_descriptor_write_writedata,
                                                reset_n,

                                               // outputs:
                                                lcd_sgdma_descriptor_write_address_to_slave,
                                                lcd_sgdma_descriptor_write_waitrequest
                                             )
;

  output  [ 31: 0] lcd_sgdma_descriptor_write_address_to_slave;
  output           lcd_sgdma_descriptor_write_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s2_end_xfer;
  input   [ 31: 0] lcd_sgdma_descriptor_write_address;
  input            lcd_sgdma_descriptor_write_granted_descriptor_memory_s2;
  input            lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2;
  input            lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;
  input            lcd_sgdma_descriptor_write_write;
  input   [ 31: 0] lcd_sgdma_descriptor_write_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 31: 0] lcd_sgdma_descriptor_write_address_last_time;
  wire    [ 31: 0] lcd_sgdma_descriptor_write_address_to_slave;
  wire             lcd_sgdma_descriptor_write_run;
  wire             lcd_sgdma_descriptor_write_waitrequest;
  reg              lcd_sgdma_descriptor_write_write_last_time;
  reg     [ 31: 0] lcd_sgdma_descriptor_write_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2 | ~lcd_sgdma_descriptor_write_requests_descriptor_memory_s2) & (lcd_sgdma_descriptor_write_granted_descriptor_memory_s2 | ~lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2) & ((~lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2 | ~(lcd_sgdma_descriptor_write_write) | (1 & (lcd_sgdma_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign lcd_sgdma_descriptor_write_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign lcd_sgdma_descriptor_write_address_to_slave = {20'b100010000000000,
    lcd_sgdma_descriptor_write_address[11 : 0]};

  //actual waitrequest port, which is an e_assign
  assign lcd_sgdma_descriptor_write_waitrequest = ~lcd_sgdma_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_sgdma_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_write_address_last_time <= 0;
      else 
        lcd_sgdma_descriptor_write_address_last_time <= lcd_sgdma_descriptor_write_address;
    end


  //lcd_sgdma/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= lcd_sgdma_descriptor_write_waitrequest & (lcd_sgdma_descriptor_write_write);
    end


  //lcd_sgdma_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_descriptor_write_address != lcd_sgdma_descriptor_write_address_last_time))
        begin
          $write("%0d ns: lcd_sgdma_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //lcd_sgdma_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_write_write_last_time <= 0;
      else 
        lcd_sgdma_descriptor_write_write_last_time <= lcd_sgdma_descriptor_write_write;
    end


  //lcd_sgdma_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_descriptor_write_write != lcd_sgdma_descriptor_write_write_last_time))
        begin
          $write("%0d ns: lcd_sgdma_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //lcd_sgdma_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_descriptor_write_writedata_last_time <= 0;
      else 
        lcd_sgdma_descriptor_write_writedata_last_time <= lcd_sgdma_descriptor_write_writedata;
    end


  //lcd_sgdma_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_descriptor_write_writedata != lcd_sgdma_descriptor_write_writedata_last_time) & lcd_sgdma_descriptor_write_write)
        begin
          $write("%0d ns: lcd_sgdma_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_sgdma_m_read_arbitrator (
                                     // inputs:
                                      clk,
                                      d1_frame_buffer_pipeline_bridge_s1_end_xfer,
                                      frame_buffer_pipeline_bridge_s1_readdata_from_sa,
                                      frame_buffer_pipeline_bridge_s1_waitrequest_from_sa,
                                      lcd_sgdma_m_read_address,
                                      lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1,
                                      lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1,
                                      lcd_sgdma_m_read_read,
                                      lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1,
                                      lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                      lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1,
                                      reset_n,

                                     // outputs:
                                      lcd_sgdma_m_read_address_to_slave,
                                      lcd_sgdma_m_read_latency_counter,
                                      lcd_sgdma_m_read_readdata,
                                      lcd_sgdma_m_read_readdatavalid,
                                      lcd_sgdma_m_read_waitrequest
                                   )
;

  output  [ 31: 0] lcd_sgdma_m_read_address_to_slave;
  output           lcd_sgdma_m_read_latency_counter;
  output  [ 31: 0] lcd_sgdma_m_read_readdata;
  output           lcd_sgdma_m_read_readdatavalid;
  output           lcd_sgdma_m_read_waitrequest;
  input            clk;
  input            d1_frame_buffer_pipeline_bridge_s1_end_xfer;
  input   [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata_from_sa;
  input            frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;
  input   [ 31: 0] lcd_sgdma_m_read_address;
  input            lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1;
  input            lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1;
  input            lcd_sgdma_m_read_read;
  input            lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1;
  input            lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  reg     [ 31: 0] lcd_sgdma_m_read_address_last_time;
  wire    [ 31: 0] lcd_sgdma_m_read_address_to_slave;
  wire             lcd_sgdma_m_read_is_granted_some_slave;
  reg              lcd_sgdma_m_read_latency_counter;
  reg              lcd_sgdma_m_read_read_but_no_slave_selected;
  reg              lcd_sgdma_m_read_read_last_time;
  wire    [ 31: 0] lcd_sgdma_m_read_readdata;
  wire             lcd_sgdma_m_read_readdatavalid;
  wire             lcd_sgdma_m_read_run;
  wire             lcd_sgdma_m_read_waitrequest;
  wire             p1_lcd_sgdma_m_read_latency_counter;
  wire             pre_flush_lcd_sgdma_m_read_readdatavalid;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1 | ~lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1) & (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1 | ~lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1) & ((~lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1 | ~(lcd_sgdma_m_read_read) | (1 & ~frame_buffer_pipeline_bridge_s1_waitrequest_from_sa & (lcd_sgdma_m_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign lcd_sgdma_m_read_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign lcd_sgdma_m_read_address_to_slave = {7'b0,
    lcd_sgdma_m_read_address[24 : 0]};

  //lcd_sgdma_m_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_m_read_read_but_no_slave_selected <= 0;
      else 
        lcd_sgdma_m_read_read_but_no_slave_selected <= lcd_sgdma_m_read_read & lcd_sgdma_m_read_run & ~lcd_sgdma_m_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign lcd_sgdma_m_read_is_granted_some_slave = lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_lcd_sgdma_m_read_readdatavalid = lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign lcd_sgdma_m_read_readdatavalid = lcd_sgdma_m_read_read_but_no_slave_selected |
    pre_flush_lcd_sgdma_m_read_readdatavalid;

  //lcd_sgdma/m_read readdata mux, which is an e_mux
  assign lcd_sgdma_m_read_readdata = frame_buffer_pipeline_bridge_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign lcd_sgdma_m_read_waitrequest = ~lcd_sgdma_m_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_m_read_latency_counter <= 0;
      else 
        lcd_sgdma_m_read_latency_counter <= p1_lcd_sgdma_m_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_lcd_sgdma_m_read_latency_counter = ((lcd_sgdma_m_read_run & lcd_sgdma_m_read_read))? latency_load_value :
    (lcd_sgdma_m_read_latency_counter)? lcd_sgdma_m_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //lcd_sgdma_m_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_m_read_address_last_time <= 0;
      else 
        lcd_sgdma_m_read_address_last_time <= lcd_sgdma_m_read_address;
    end


  //lcd_sgdma/m_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= lcd_sgdma_m_read_waitrequest & (lcd_sgdma_m_read_read);
    end


  //lcd_sgdma_m_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_m_read_address != lcd_sgdma_m_read_address_last_time))
        begin
          $write("%0d ns: lcd_sgdma_m_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //lcd_sgdma_m_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          lcd_sgdma_m_read_read_last_time <= 0;
      else 
        lcd_sgdma_m_read_read_last_time <= lcd_sgdma_m_read_read;
    end


  //lcd_sgdma_m_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (lcd_sgdma_m_read_read != lcd_sgdma_m_read_read_last_time))
        begin
          $write("%0d ns: lcd_sgdma_m_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_sgdma_out_arbitrator (
                                  // inputs:
                                   clk,
                                   lcd_pixel_converter_in_ready_from_sa,
                                   lcd_sgdma_out_data,
                                   lcd_sgdma_out_empty,
                                   lcd_sgdma_out_endofpacket,
                                   lcd_sgdma_out_startofpacket,
                                   lcd_sgdma_out_valid,
                                   reset_n,

                                  // outputs:
                                   lcd_sgdma_out_ready
                                )
;

  output           lcd_sgdma_out_ready;
  input            clk;
  input            lcd_pixel_converter_in_ready_from_sa;
  input   [ 31: 0] lcd_sgdma_out_data;
  input   [  1: 0] lcd_sgdma_out_empty;
  input            lcd_sgdma_out_endofpacket;
  input            lcd_sgdma_out_startofpacket;
  input            lcd_sgdma_out_valid;
  input            reset_n;

  wire             lcd_sgdma_out_ready;
  //mux lcd_sgdma_out_ready, which is an e_mux
  assign lcd_sgdma_out_ready = lcd_pixel_converter_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_ta_fifo_to_sequencer_in_arbitrator (
                                                // inputs:
                                                 clk,
                                                 lcd_on_chip_memory_fifo_out_data,
                                                 lcd_on_chip_memory_fifo_out_endofpacket,
                                                 lcd_on_chip_memory_fifo_out_startofpacket,
                                                 lcd_on_chip_memory_fifo_out_valid,
                                                 lcd_ta_fifo_to_sequencer_in_ready,
                                                 reset_n,

                                                // outputs:
                                                 lcd_ta_fifo_to_sequencer_in_data,
                                                 lcd_ta_fifo_to_sequencer_in_endofpacket,
                                                 lcd_ta_fifo_to_sequencer_in_ready_from_sa,
                                                 lcd_ta_fifo_to_sequencer_in_reset_n,
                                                 lcd_ta_fifo_to_sequencer_in_startofpacket,
                                                 lcd_ta_fifo_to_sequencer_in_valid
                                              )
;

  output  [  7: 0] lcd_ta_fifo_to_sequencer_in_data;
  output           lcd_ta_fifo_to_sequencer_in_endofpacket;
  output           lcd_ta_fifo_to_sequencer_in_ready_from_sa;
  output           lcd_ta_fifo_to_sequencer_in_reset_n;
  output           lcd_ta_fifo_to_sequencer_in_startofpacket;
  output           lcd_ta_fifo_to_sequencer_in_valid;
  input            clk;
  input   [  7: 0] lcd_on_chip_memory_fifo_out_data;
  input            lcd_on_chip_memory_fifo_out_endofpacket;
  input            lcd_on_chip_memory_fifo_out_startofpacket;
  input            lcd_on_chip_memory_fifo_out_valid;
  input            lcd_ta_fifo_to_sequencer_in_ready;
  input            reset_n;

  wire    [  7: 0] lcd_ta_fifo_to_sequencer_in_data;
  wire             lcd_ta_fifo_to_sequencer_in_endofpacket;
  wire             lcd_ta_fifo_to_sequencer_in_ready_from_sa;
  wire             lcd_ta_fifo_to_sequencer_in_reset_n;
  wire             lcd_ta_fifo_to_sequencer_in_startofpacket;
  wire             lcd_ta_fifo_to_sequencer_in_valid;
  //mux lcd_ta_fifo_to_sequencer_in_data, which is an e_mux
  assign lcd_ta_fifo_to_sequencer_in_data = lcd_on_chip_memory_fifo_out_data;

  //mux lcd_ta_fifo_to_sequencer_in_endofpacket, which is an e_mux
  assign lcd_ta_fifo_to_sequencer_in_endofpacket = lcd_on_chip_memory_fifo_out_endofpacket;

  //assign lcd_ta_fifo_to_sequencer_in_ready_from_sa = lcd_ta_fifo_to_sequencer_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_ta_fifo_to_sequencer_in_ready_from_sa = lcd_ta_fifo_to_sequencer_in_ready;

  //mux lcd_ta_fifo_to_sequencer_in_startofpacket, which is an e_mux
  assign lcd_ta_fifo_to_sequencer_in_startofpacket = lcd_on_chip_memory_fifo_out_startofpacket;

  //mux lcd_ta_fifo_to_sequencer_in_valid, which is an e_mux
  assign lcd_ta_fifo_to_sequencer_in_valid = lcd_on_chip_memory_fifo_out_valid;

  //lcd_ta_fifo_to_sequencer_in_reset_n assignment, which is an e_assign
  assign lcd_ta_fifo_to_sequencer_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_ta_fifo_to_sequencer_out_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  lcd_data_format_adapter_1_in_ready_from_sa,
                                                  lcd_ta_fifo_to_sequencer_out_data,
                                                  lcd_ta_fifo_to_sequencer_out_endofpacket,
                                                  lcd_ta_fifo_to_sequencer_out_startofpacket,
                                                  lcd_ta_fifo_to_sequencer_out_valid,
                                                  reset_n,

                                                 // outputs:
                                                  lcd_ta_fifo_to_sequencer_out_ready
                                               )
;

  output           lcd_ta_fifo_to_sequencer_out_ready;
  input            clk;
  input            lcd_data_format_adapter_1_in_ready_from_sa;
  input   [  7: 0] lcd_ta_fifo_to_sequencer_out_data;
  input            lcd_ta_fifo_to_sequencer_out_endofpacket;
  input            lcd_ta_fifo_to_sequencer_out_startofpacket;
  input            lcd_ta_fifo_to_sequencer_out_valid;
  input            reset_n;

  wire             lcd_ta_fifo_to_sequencer_out_ready;
  //mux lcd_ta_fifo_to_sequencer_out_ready, which is an e_mux
  assign lcd_ta_fifo_to_sequencer_out_ready = lcd_data_format_adapter_1_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_ta_formatter_to_fifo_in_arbitrator (
                                                // inputs:
                                                 clk,
                                                 lcd_data_format_adapter_out_data,
                                                 lcd_data_format_adapter_out_endofpacket,
                                                 lcd_data_format_adapter_out_startofpacket,
                                                 lcd_data_format_adapter_out_valid,
                                                 lcd_ta_formatter_to_fifo_in_ready,
                                                 reset_n,

                                                // outputs:
                                                 lcd_ta_formatter_to_fifo_in_data,
                                                 lcd_ta_formatter_to_fifo_in_endofpacket,
                                                 lcd_ta_formatter_to_fifo_in_ready_from_sa,
                                                 lcd_ta_formatter_to_fifo_in_reset_n,
                                                 lcd_ta_formatter_to_fifo_in_startofpacket,
                                                 lcd_ta_formatter_to_fifo_in_valid
                                              )
;

  output  [  7: 0] lcd_ta_formatter_to_fifo_in_data;
  output           lcd_ta_formatter_to_fifo_in_endofpacket;
  output           lcd_ta_formatter_to_fifo_in_ready_from_sa;
  output           lcd_ta_formatter_to_fifo_in_reset_n;
  output           lcd_ta_formatter_to_fifo_in_startofpacket;
  output           lcd_ta_formatter_to_fifo_in_valid;
  input            clk;
  input   [  7: 0] lcd_data_format_adapter_out_data;
  input            lcd_data_format_adapter_out_endofpacket;
  input            lcd_data_format_adapter_out_startofpacket;
  input            lcd_data_format_adapter_out_valid;
  input            lcd_ta_formatter_to_fifo_in_ready;
  input            reset_n;

  wire    [  7: 0] lcd_ta_formatter_to_fifo_in_data;
  wire             lcd_ta_formatter_to_fifo_in_endofpacket;
  wire             lcd_ta_formatter_to_fifo_in_ready_from_sa;
  wire             lcd_ta_formatter_to_fifo_in_reset_n;
  wire             lcd_ta_formatter_to_fifo_in_startofpacket;
  wire             lcd_ta_formatter_to_fifo_in_valid;
  //mux lcd_ta_formatter_to_fifo_in_data, which is an e_mux
  assign lcd_ta_formatter_to_fifo_in_data = lcd_data_format_adapter_out_data;

  //mux lcd_ta_formatter_to_fifo_in_endofpacket, which is an e_mux
  assign lcd_ta_formatter_to_fifo_in_endofpacket = lcd_data_format_adapter_out_endofpacket;

  //assign lcd_ta_formatter_to_fifo_in_ready_from_sa = lcd_ta_formatter_to_fifo_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_ta_formatter_to_fifo_in_ready_from_sa = lcd_ta_formatter_to_fifo_in_ready;

  //mux lcd_ta_formatter_to_fifo_in_startofpacket, which is an e_mux
  assign lcd_ta_formatter_to_fifo_in_startofpacket = lcd_data_format_adapter_out_startofpacket;

  //mux lcd_ta_formatter_to_fifo_in_valid, which is an e_mux
  assign lcd_ta_formatter_to_fifo_in_valid = lcd_data_format_adapter_out_valid;

  //lcd_ta_formatter_to_fifo_in_reset_n assignment, which is an e_assign
  assign lcd_ta_formatter_to_fifo_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_ta_formatter_to_fifo_out_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  lcd_on_chip_memory_fifo_in_ready_from_sa,
                                                  lcd_ta_formatter_to_fifo_out_data,
                                                  lcd_ta_formatter_to_fifo_out_endofpacket,
                                                  lcd_ta_formatter_to_fifo_out_startofpacket,
                                                  lcd_ta_formatter_to_fifo_out_valid,
                                                  reset_n,

                                                 // outputs:
                                                  lcd_ta_formatter_to_fifo_out_ready
                                               )
;

  output           lcd_ta_formatter_to_fifo_out_ready;
  input            clk;
  input            lcd_on_chip_memory_fifo_in_ready_from_sa;
  input   [  7: 0] lcd_ta_formatter_to_fifo_out_data;
  input            lcd_ta_formatter_to_fifo_out_endofpacket;
  input            lcd_ta_formatter_to_fifo_out_startofpacket;
  input            lcd_ta_formatter_to_fifo_out_valid;
  input            reset_n;

  wire             lcd_ta_formatter_to_fifo_out_ready;
  //mux lcd_ta_formatter_to_fifo_out_ready, which is an e_mux
  assign lcd_ta_formatter_to_fifo_out_ready = lcd_on_chip_memory_fifo_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lcd_video_sequencer_in_arbitrator (
                                           // inputs:
                                            clk,
                                            lcd_data_format_adapter_1_out_data,
                                            lcd_data_format_adapter_1_out_empty,
                                            lcd_data_format_adapter_1_out_endofpacket,
                                            lcd_data_format_adapter_1_out_startofpacket,
                                            lcd_data_format_adapter_1_out_valid,
                                            lcd_video_sequencer_in_ready,
                                            reset_n,

                                           // outputs:
                                            lcd_video_sequencer_in_data,
                                            lcd_video_sequencer_in_empty,
                                            lcd_video_sequencer_in_endofpacket,
                                            lcd_video_sequencer_in_ready_from_sa,
                                            lcd_video_sequencer_in_reset_n,
                                            lcd_video_sequencer_in_startofpacket,
                                            lcd_video_sequencer_in_valid
                                         )
;

  output  [  7: 0] lcd_video_sequencer_in_data;
  output           lcd_video_sequencer_in_empty;
  output           lcd_video_sequencer_in_endofpacket;
  output           lcd_video_sequencer_in_ready_from_sa;
  output           lcd_video_sequencer_in_reset_n;
  output           lcd_video_sequencer_in_startofpacket;
  output           lcd_video_sequencer_in_valid;
  input            clk;
  input   [  7: 0] lcd_data_format_adapter_1_out_data;
  input            lcd_data_format_adapter_1_out_empty;
  input            lcd_data_format_adapter_1_out_endofpacket;
  input            lcd_data_format_adapter_1_out_startofpacket;
  input            lcd_data_format_adapter_1_out_valid;
  input            lcd_video_sequencer_in_ready;
  input            reset_n;

  wire    [  7: 0] lcd_video_sequencer_in_data;
  wire             lcd_video_sequencer_in_empty;
  wire             lcd_video_sequencer_in_endofpacket;
  wire             lcd_video_sequencer_in_ready_from_sa;
  wire             lcd_video_sequencer_in_reset_n;
  wire             lcd_video_sequencer_in_startofpacket;
  wire             lcd_video_sequencer_in_valid;
  //mux lcd_video_sequencer_in_data, which is an e_mux
  assign lcd_video_sequencer_in_data = lcd_data_format_adapter_1_out_data;

  //mux lcd_video_sequencer_in_empty, which is an e_mux
  assign lcd_video_sequencer_in_empty = lcd_data_format_adapter_1_out_empty;

  //mux lcd_video_sequencer_in_endofpacket, which is an e_mux
  assign lcd_video_sequencer_in_endofpacket = lcd_data_format_adapter_1_out_endofpacket;

  //assign lcd_video_sequencer_in_ready_from_sa = lcd_video_sequencer_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign lcd_video_sequencer_in_ready_from_sa = lcd_video_sequencer_in_ready;

  //mux lcd_video_sequencer_in_startofpacket, which is an e_mux
  assign lcd_video_sequencer_in_startofpacket = lcd_data_format_adapter_1_out_startofpacket;

  //mux lcd_video_sequencer_in_valid, which is an e_mux
  assign lcd_video_sequencer_in_valid = lcd_data_format_adapter_1_out_valid;

  //lcd_video_sequencer_in_reset_n assignment, which is an e_assign
  assign lcd_video_sequencer_in_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pio_id_eeprom_dat_s1_arbitrator (
                                         // inputs:
                                          clk,
                                          clock_crossing_bridge_m1_address_to_slave,
                                          clock_crossing_bridge_m1_latency_counter,
                                          clock_crossing_bridge_m1_nativeaddress,
                                          clock_crossing_bridge_m1_read,
                                          clock_crossing_bridge_m1_write,
                                          clock_crossing_bridge_m1_writedata,
                                          pio_id_eeprom_dat_s1_readdata,
                                          reset_n,

                                         // outputs:
                                          clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1,
                                          clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1,
                                          clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1,
                                          clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1,
                                          d1_pio_id_eeprom_dat_s1_end_xfer,
                                          pio_id_eeprom_dat_s1_address,
                                          pio_id_eeprom_dat_s1_chipselect,
                                          pio_id_eeprom_dat_s1_readdata_from_sa,
                                          pio_id_eeprom_dat_s1_reset_n,
                                          pio_id_eeprom_dat_s1_write_n,
                                          pio_id_eeprom_dat_s1_writedata
                                       )
;

  output           clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1;
  output           clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1;
  output           clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1;
  output           clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1;
  output           d1_pio_id_eeprom_dat_s1_end_xfer;
  output  [  1: 0] pio_id_eeprom_dat_s1_address;
  output           pio_id_eeprom_dat_s1_chipselect;
  output  [ 31: 0] pio_id_eeprom_dat_s1_readdata_from_sa;
  output           pio_id_eeprom_dat_s1_reset_n;
  output           pio_id_eeprom_dat_s1_write_n;
  output  [ 31: 0] pio_id_eeprom_dat_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] pio_id_eeprom_dat_s1_readdata;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_saved_grant_pio_id_eeprom_dat_s1;
  reg              d1_pio_id_eeprom_dat_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] pio_id_eeprom_dat_s1_address;
  wire             pio_id_eeprom_dat_s1_allgrants;
  wire             pio_id_eeprom_dat_s1_allow_new_arb_cycle;
  wire             pio_id_eeprom_dat_s1_any_bursting_master_saved_grant;
  wire             pio_id_eeprom_dat_s1_any_continuerequest;
  wire             pio_id_eeprom_dat_s1_arb_counter_enable;
  reg              pio_id_eeprom_dat_s1_arb_share_counter;
  wire             pio_id_eeprom_dat_s1_arb_share_counter_next_value;
  wire             pio_id_eeprom_dat_s1_arb_share_set_values;
  wire             pio_id_eeprom_dat_s1_beginbursttransfer_internal;
  wire             pio_id_eeprom_dat_s1_begins_xfer;
  wire             pio_id_eeprom_dat_s1_chipselect;
  wire             pio_id_eeprom_dat_s1_end_xfer;
  wire             pio_id_eeprom_dat_s1_firsttransfer;
  wire             pio_id_eeprom_dat_s1_grant_vector;
  wire             pio_id_eeprom_dat_s1_in_a_read_cycle;
  wire             pio_id_eeprom_dat_s1_in_a_write_cycle;
  wire             pio_id_eeprom_dat_s1_master_qreq_vector;
  wire             pio_id_eeprom_dat_s1_non_bursting_master_requests;
  wire    [ 31: 0] pio_id_eeprom_dat_s1_readdata_from_sa;
  reg              pio_id_eeprom_dat_s1_reg_firsttransfer;
  wire             pio_id_eeprom_dat_s1_reset_n;
  reg              pio_id_eeprom_dat_s1_slavearbiterlockenable;
  wire             pio_id_eeprom_dat_s1_slavearbiterlockenable2;
  wire             pio_id_eeprom_dat_s1_unreg_firsttransfer;
  wire             pio_id_eeprom_dat_s1_waits_for_read;
  wire             pio_id_eeprom_dat_s1_waits_for_write;
  wire             pio_id_eeprom_dat_s1_write_n;
  wire    [ 31: 0] pio_id_eeprom_dat_s1_writedata;
  wire             wait_for_pio_id_eeprom_dat_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pio_id_eeprom_dat_s1_end_xfer;
    end


  assign pio_id_eeprom_dat_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1));
  //assign pio_id_eeprom_dat_s1_readdata_from_sa = pio_id_eeprom_dat_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pio_id_eeprom_dat_s1_readdata_from_sa = pio_id_eeprom_dat_s1_readdata;

  assign clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h480) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //pio_id_eeprom_dat_s1_arb_share_counter set values, which is an e_mux
  assign pio_id_eeprom_dat_s1_arb_share_set_values = 1;

  //pio_id_eeprom_dat_s1_non_bursting_master_requests mux, which is an e_mux
  assign pio_id_eeprom_dat_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1;

  //pio_id_eeprom_dat_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pio_id_eeprom_dat_s1_any_bursting_master_saved_grant = 0;

  //pio_id_eeprom_dat_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pio_id_eeprom_dat_s1_arb_share_counter_next_value = pio_id_eeprom_dat_s1_firsttransfer ? (pio_id_eeprom_dat_s1_arb_share_set_values - 1) : |pio_id_eeprom_dat_s1_arb_share_counter ? (pio_id_eeprom_dat_s1_arb_share_counter - 1) : 0;

  //pio_id_eeprom_dat_s1_allgrants all slave grants, which is an e_mux
  assign pio_id_eeprom_dat_s1_allgrants = |pio_id_eeprom_dat_s1_grant_vector;

  //pio_id_eeprom_dat_s1_end_xfer assignment, which is an e_assign
  assign pio_id_eeprom_dat_s1_end_xfer = ~(pio_id_eeprom_dat_s1_waits_for_read | pio_id_eeprom_dat_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1 = pio_id_eeprom_dat_s1_end_xfer & (~pio_id_eeprom_dat_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pio_id_eeprom_dat_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pio_id_eeprom_dat_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1 & pio_id_eeprom_dat_s1_allgrants) | (end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1 & ~pio_id_eeprom_dat_s1_non_bursting_master_requests);

  //pio_id_eeprom_dat_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pio_id_eeprom_dat_s1_arb_share_counter <= 0;
      else if (pio_id_eeprom_dat_s1_arb_counter_enable)
          pio_id_eeprom_dat_s1_arb_share_counter <= pio_id_eeprom_dat_s1_arb_share_counter_next_value;
    end


  //pio_id_eeprom_dat_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pio_id_eeprom_dat_s1_slavearbiterlockenable <= 0;
      else if ((|pio_id_eeprom_dat_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1) | (end_xfer_arb_share_counter_term_pio_id_eeprom_dat_s1 & ~pio_id_eeprom_dat_s1_non_bursting_master_requests))
          pio_id_eeprom_dat_s1_slavearbiterlockenable <= |pio_id_eeprom_dat_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 pio_id_eeprom_dat/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = pio_id_eeprom_dat_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //pio_id_eeprom_dat_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pio_id_eeprom_dat_s1_slavearbiterlockenable2 = |pio_id_eeprom_dat_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 pio_id_eeprom_dat/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = pio_id_eeprom_dat_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //pio_id_eeprom_dat_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pio_id_eeprom_dat_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1 = clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1 = clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1 & clock_crossing_bridge_m1_read & ~pio_id_eeprom_dat_s1_waits_for_read;

  //pio_id_eeprom_dat_s1_writedata mux, which is an e_mux
  assign pio_id_eeprom_dat_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1 = clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1;

  //clock_crossing_bridge/m1 saved-grant pio_id_eeprom_dat/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_pio_id_eeprom_dat_s1 = clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1;

  //allow new arb cycle for pio_id_eeprom_dat/s1, which is an e_assign
  assign pio_id_eeprom_dat_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pio_id_eeprom_dat_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pio_id_eeprom_dat_s1_master_qreq_vector = 1;

  //pio_id_eeprom_dat_s1_reset_n assignment, which is an e_assign
  assign pio_id_eeprom_dat_s1_reset_n = reset_n;

  assign pio_id_eeprom_dat_s1_chipselect = clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1;
  //pio_id_eeprom_dat_s1_firsttransfer first transaction, which is an e_assign
  assign pio_id_eeprom_dat_s1_firsttransfer = pio_id_eeprom_dat_s1_begins_xfer ? pio_id_eeprom_dat_s1_unreg_firsttransfer : pio_id_eeprom_dat_s1_reg_firsttransfer;

  //pio_id_eeprom_dat_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pio_id_eeprom_dat_s1_unreg_firsttransfer = ~(pio_id_eeprom_dat_s1_slavearbiterlockenable & pio_id_eeprom_dat_s1_any_continuerequest);

  //pio_id_eeprom_dat_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pio_id_eeprom_dat_s1_reg_firsttransfer <= 1'b1;
      else if (pio_id_eeprom_dat_s1_begins_xfer)
          pio_id_eeprom_dat_s1_reg_firsttransfer <= pio_id_eeprom_dat_s1_unreg_firsttransfer;
    end


  //pio_id_eeprom_dat_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pio_id_eeprom_dat_s1_beginbursttransfer_internal = pio_id_eeprom_dat_s1_begins_xfer;

  //~pio_id_eeprom_dat_s1_write_n assignment, which is an e_mux
  assign pio_id_eeprom_dat_s1_write_n = ~(clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1 & clock_crossing_bridge_m1_write);

  //pio_id_eeprom_dat_s1_address mux, which is an e_mux
  assign pio_id_eeprom_dat_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_pio_id_eeprom_dat_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pio_id_eeprom_dat_s1_end_xfer <= 1;
      else 
        d1_pio_id_eeprom_dat_s1_end_xfer <= pio_id_eeprom_dat_s1_end_xfer;
    end


  //pio_id_eeprom_dat_s1_waits_for_read in a cycle, which is an e_mux
  assign pio_id_eeprom_dat_s1_waits_for_read = pio_id_eeprom_dat_s1_in_a_read_cycle & pio_id_eeprom_dat_s1_begins_xfer;

  //pio_id_eeprom_dat_s1_in_a_read_cycle assignment, which is an e_assign
  assign pio_id_eeprom_dat_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pio_id_eeprom_dat_s1_in_a_read_cycle;

  //pio_id_eeprom_dat_s1_waits_for_write in a cycle, which is an e_mux
  assign pio_id_eeprom_dat_s1_waits_for_write = pio_id_eeprom_dat_s1_in_a_write_cycle & 0;

  //pio_id_eeprom_dat_s1_in_a_write_cycle assignment, which is an e_assign
  assign pio_id_eeprom_dat_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pio_id_eeprom_dat_s1_in_a_write_cycle;

  assign wait_for_pio_id_eeprom_dat_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pio_id_eeprom_dat/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pio_id_eeprom_scl_s1_arbitrator (
                                         // inputs:
                                          clk,
                                          clock_crossing_bridge_m1_address_to_slave,
                                          clock_crossing_bridge_m1_latency_counter,
                                          clock_crossing_bridge_m1_nativeaddress,
                                          clock_crossing_bridge_m1_read,
                                          clock_crossing_bridge_m1_write,
                                          clock_crossing_bridge_m1_writedata,
                                          pio_id_eeprom_scl_s1_readdata,
                                          reset_n,

                                         // outputs:
                                          clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1,
                                          clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1,
                                          clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1,
                                          clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1,
                                          d1_pio_id_eeprom_scl_s1_end_xfer,
                                          pio_id_eeprom_scl_s1_address,
                                          pio_id_eeprom_scl_s1_chipselect,
                                          pio_id_eeprom_scl_s1_readdata_from_sa,
                                          pio_id_eeprom_scl_s1_reset_n,
                                          pio_id_eeprom_scl_s1_write_n,
                                          pio_id_eeprom_scl_s1_writedata
                                       )
;

  output           clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1;
  output           clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1;
  output           clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1;
  output           clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1;
  output           d1_pio_id_eeprom_scl_s1_end_xfer;
  output  [  1: 0] pio_id_eeprom_scl_s1_address;
  output           pio_id_eeprom_scl_s1_chipselect;
  output  [ 31: 0] pio_id_eeprom_scl_s1_readdata_from_sa;
  output           pio_id_eeprom_scl_s1_reset_n;
  output           pio_id_eeprom_scl_s1_write_n;
  output  [ 31: 0] pio_id_eeprom_scl_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input   [ 31: 0] pio_id_eeprom_scl_s1_readdata;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_saved_grant_pio_id_eeprom_scl_s1;
  reg              d1_pio_id_eeprom_scl_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] pio_id_eeprom_scl_s1_address;
  wire             pio_id_eeprom_scl_s1_allgrants;
  wire             pio_id_eeprom_scl_s1_allow_new_arb_cycle;
  wire             pio_id_eeprom_scl_s1_any_bursting_master_saved_grant;
  wire             pio_id_eeprom_scl_s1_any_continuerequest;
  wire             pio_id_eeprom_scl_s1_arb_counter_enable;
  reg              pio_id_eeprom_scl_s1_arb_share_counter;
  wire             pio_id_eeprom_scl_s1_arb_share_counter_next_value;
  wire             pio_id_eeprom_scl_s1_arb_share_set_values;
  wire             pio_id_eeprom_scl_s1_beginbursttransfer_internal;
  wire             pio_id_eeprom_scl_s1_begins_xfer;
  wire             pio_id_eeprom_scl_s1_chipselect;
  wire             pio_id_eeprom_scl_s1_end_xfer;
  wire             pio_id_eeprom_scl_s1_firsttransfer;
  wire             pio_id_eeprom_scl_s1_grant_vector;
  wire             pio_id_eeprom_scl_s1_in_a_read_cycle;
  wire             pio_id_eeprom_scl_s1_in_a_write_cycle;
  wire             pio_id_eeprom_scl_s1_master_qreq_vector;
  wire             pio_id_eeprom_scl_s1_non_bursting_master_requests;
  wire    [ 31: 0] pio_id_eeprom_scl_s1_readdata_from_sa;
  reg              pio_id_eeprom_scl_s1_reg_firsttransfer;
  wire             pio_id_eeprom_scl_s1_reset_n;
  reg              pio_id_eeprom_scl_s1_slavearbiterlockenable;
  wire             pio_id_eeprom_scl_s1_slavearbiterlockenable2;
  wire             pio_id_eeprom_scl_s1_unreg_firsttransfer;
  wire             pio_id_eeprom_scl_s1_waits_for_read;
  wire             pio_id_eeprom_scl_s1_waits_for_write;
  wire             pio_id_eeprom_scl_s1_write_n;
  wire    [ 31: 0] pio_id_eeprom_scl_s1_writedata;
  wire             wait_for_pio_id_eeprom_scl_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pio_id_eeprom_scl_s1_end_xfer;
    end


  assign pio_id_eeprom_scl_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1));
  //assign pio_id_eeprom_scl_s1_readdata_from_sa = pio_id_eeprom_scl_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pio_id_eeprom_scl_s1_readdata_from_sa = pio_id_eeprom_scl_s1_readdata;

  assign clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h500) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //pio_id_eeprom_scl_s1_arb_share_counter set values, which is an e_mux
  assign pio_id_eeprom_scl_s1_arb_share_set_values = 1;

  //pio_id_eeprom_scl_s1_non_bursting_master_requests mux, which is an e_mux
  assign pio_id_eeprom_scl_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1;

  //pio_id_eeprom_scl_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pio_id_eeprom_scl_s1_any_bursting_master_saved_grant = 0;

  //pio_id_eeprom_scl_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pio_id_eeprom_scl_s1_arb_share_counter_next_value = pio_id_eeprom_scl_s1_firsttransfer ? (pio_id_eeprom_scl_s1_arb_share_set_values - 1) : |pio_id_eeprom_scl_s1_arb_share_counter ? (pio_id_eeprom_scl_s1_arb_share_counter - 1) : 0;

  //pio_id_eeprom_scl_s1_allgrants all slave grants, which is an e_mux
  assign pio_id_eeprom_scl_s1_allgrants = |pio_id_eeprom_scl_s1_grant_vector;

  //pio_id_eeprom_scl_s1_end_xfer assignment, which is an e_assign
  assign pio_id_eeprom_scl_s1_end_xfer = ~(pio_id_eeprom_scl_s1_waits_for_read | pio_id_eeprom_scl_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1 = pio_id_eeprom_scl_s1_end_xfer & (~pio_id_eeprom_scl_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pio_id_eeprom_scl_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pio_id_eeprom_scl_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1 & pio_id_eeprom_scl_s1_allgrants) | (end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1 & ~pio_id_eeprom_scl_s1_non_bursting_master_requests);

  //pio_id_eeprom_scl_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pio_id_eeprom_scl_s1_arb_share_counter <= 0;
      else if (pio_id_eeprom_scl_s1_arb_counter_enable)
          pio_id_eeprom_scl_s1_arb_share_counter <= pio_id_eeprom_scl_s1_arb_share_counter_next_value;
    end


  //pio_id_eeprom_scl_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pio_id_eeprom_scl_s1_slavearbiterlockenable <= 0;
      else if ((|pio_id_eeprom_scl_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1) | (end_xfer_arb_share_counter_term_pio_id_eeprom_scl_s1 & ~pio_id_eeprom_scl_s1_non_bursting_master_requests))
          pio_id_eeprom_scl_s1_slavearbiterlockenable <= |pio_id_eeprom_scl_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 pio_id_eeprom_scl/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = pio_id_eeprom_scl_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //pio_id_eeprom_scl_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pio_id_eeprom_scl_s1_slavearbiterlockenable2 = |pio_id_eeprom_scl_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 pio_id_eeprom_scl/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = pio_id_eeprom_scl_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //pio_id_eeprom_scl_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pio_id_eeprom_scl_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1 = clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1 = clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1 & clock_crossing_bridge_m1_read & ~pio_id_eeprom_scl_s1_waits_for_read;

  //pio_id_eeprom_scl_s1_writedata mux, which is an e_mux
  assign pio_id_eeprom_scl_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1 = clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1;

  //clock_crossing_bridge/m1 saved-grant pio_id_eeprom_scl/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_pio_id_eeprom_scl_s1 = clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1;

  //allow new arb cycle for pio_id_eeprom_scl/s1, which is an e_assign
  assign pio_id_eeprom_scl_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pio_id_eeprom_scl_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pio_id_eeprom_scl_s1_master_qreq_vector = 1;

  //pio_id_eeprom_scl_s1_reset_n assignment, which is an e_assign
  assign pio_id_eeprom_scl_s1_reset_n = reset_n;

  assign pio_id_eeprom_scl_s1_chipselect = clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1;
  //pio_id_eeprom_scl_s1_firsttransfer first transaction, which is an e_assign
  assign pio_id_eeprom_scl_s1_firsttransfer = pio_id_eeprom_scl_s1_begins_xfer ? pio_id_eeprom_scl_s1_unreg_firsttransfer : pio_id_eeprom_scl_s1_reg_firsttransfer;

  //pio_id_eeprom_scl_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pio_id_eeprom_scl_s1_unreg_firsttransfer = ~(pio_id_eeprom_scl_s1_slavearbiterlockenable & pio_id_eeprom_scl_s1_any_continuerequest);

  //pio_id_eeprom_scl_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pio_id_eeprom_scl_s1_reg_firsttransfer <= 1'b1;
      else if (pio_id_eeprom_scl_s1_begins_xfer)
          pio_id_eeprom_scl_s1_reg_firsttransfer <= pio_id_eeprom_scl_s1_unreg_firsttransfer;
    end


  //pio_id_eeprom_scl_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pio_id_eeprom_scl_s1_beginbursttransfer_internal = pio_id_eeprom_scl_s1_begins_xfer;

  //~pio_id_eeprom_scl_s1_write_n assignment, which is an e_mux
  assign pio_id_eeprom_scl_s1_write_n = ~(clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1 & clock_crossing_bridge_m1_write);

  //pio_id_eeprom_scl_s1_address mux, which is an e_mux
  assign pio_id_eeprom_scl_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_pio_id_eeprom_scl_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pio_id_eeprom_scl_s1_end_xfer <= 1;
      else 
        d1_pio_id_eeprom_scl_s1_end_xfer <= pio_id_eeprom_scl_s1_end_xfer;
    end


  //pio_id_eeprom_scl_s1_waits_for_read in a cycle, which is an e_mux
  assign pio_id_eeprom_scl_s1_waits_for_read = pio_id_eeprom_scl_s1_in_a_read_cycle & pio_id_eeprom_scl_s1_begins_xfer;

  //pio_id_eeprom_scl_s1_in_a_read_cycle assignment, which is an e_assign
  assign pio_id_eeprom_scl_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pio_id_eeprom_scl_s1_in_a_read_cycle;

  //pio_id_eeprom_scl_s1_waits_for_write in a cycle, which is an e_mux
  assign pio_id_eeprom_scl_s1_waits_for_write = pio_id_eeprom_scl_s1_in_a_write_cycle & 0;

  //pio_id_eeprom_scl_s1_in_a_write_cycle assignment, which is an e_assign
  assign pio_id_eeprom_scl_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pio_id_eeprom_scl_s1_in_a_write_cycle;

  assign wait_for_pio_id_eeprom_scl_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pio_id_eeprom_scl/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  wire             full_54;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_53;
  assign empty = !full_0;
  assign full_54 = 0;
  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    0;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  reg              full_48;
  reg              full_49;
  reg              full_5;
  reg              full_50;
  reg              full_51;
  reg              full_52;
  reg              full_53;
  wire             full_54;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p48_full_48;
  wire             p48_stage_48;
  wire             p49_full_49;
  wire             p49_stage_49;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p50_full_50;
  wire             p50_stage_50;
  wire             p51_full_51;
  wire             p51_stage_51;
  wire             p52_full_52;
  wire             p52_stage_52;
  wire             p53_full_53;
  wire             p53_stage_53;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_48;
  reg              stage_49;
  reg              stage_5;
  reg              stage_50;
  reg              stage_51;
  reg              stage_52;
  reg              stage_53;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_53;
  assign empty = !full_0;
  assign full_54 = 0;
  //data_53, which is an e_mux
  assign p53_stage_53 = ((full_54 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_53 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_53))
          if (sync_reset & full_53 & !((full_54 == 0) & read & write))
              stage_53 <= 0;
          else 
            stage_53 <= p53_stage_53;
    end


  //control_53, which is an e_mux
  assign p53_full_53 = ((read & !write) == 0)? full_52 :
    0;

  //control_reg_53, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_53 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_53 <= 0;
          else 
            full_53 <= p53_full_53;
    end


  //data_52, which is an e_mux
  assign p52_stage_52 = ((full_53 & ~clear_fifo) == 0)? data_in :
    stage_53;

  //data_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_52 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_52))
          if (sync_reset & full_52 & !((full_53 == 0) & read & write))
              stage_52 <= 0;
          else 
            stage_52 <= p52_stage_52;
    end


  //control_52, which is an e_mux
  assign p52_full_52 = ((read & !write) == 0)? full_51 :
    full_53;

  //control_reg_52, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_52 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_52 <= 0;
          else 
            full_52 <= p52_full_52;
    end


  //data_51, which is an e_mux
  assign p51_stage_51 = ((full_52 & ~clear_fifo) == 0)? data_in :
    stage_52;

  //data_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_51 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_51))
          if (sync_reset & full_51 & !((full_52 == 0) & read & write))
              stage_51 <= 0;
          else 
            stage_51 <= p51_stage_51;
    end


  //control_51, which is an e_mux
  assign p51_full_51 = ((read & !write) == 0)? full_50 :
    full_52;

  //control_reg_51, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_51 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_51 <= 0;
          else 
            full_51 <= p51_full_51;
    end


  //data_50, which is an e_mux
  assign p50_stage_50 = ((full_51 & ~clear_fifo) == 0)? data_in :
    stage_51;

  //data_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_50 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_50))
          if (sync_reset & full_50 & !((full_51 == 0) & read & write))
              stage_50 <= 0;
          else 
            stage_50 <= p50_stage_50;
    end


  //control_50, which is an e_mux
  assign p50_full_50 = ((read & !write) == 0)? full_49 :
    full_51;

  //control_reg_50, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_50 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_50 <= 0;
          else 
            full_50 <= p50_full_50;
    end


  //data_49, which is an e_mux
  assign p49_stage_49 = ((full_50 & ~clear_fifo) == 0)? data_in :
    stage_50;

  //data_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_49 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_49))
          if (sync_reset & full_49 & !((full_50 == 0) & read & write))
              stage_49 <= 0;
          else 
            stage_49 <= p49_stage_49;
    end


  //control_49, which is an e_mux
  assign p49_full_49 = ((read & !write) == 0)? full_48 :
    full_50;

  //control_reg_49, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_49 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_49 <= 0;
          else 
            full_49 <= p49_full_49;
    end


  //data_48, which is an e_mux
  assign p48_stage_48 = ((full_49 & ~clear_fifo) == 0)? data_in :
    stage_49;

  //data_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_48 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_48))
          if (sync_reset & full_48 & !((full_49 == 0) & read & write))
              stage_48 <= 0;
          else 
            stage_48 <= p48_stage_48;
    end


  //control_48, which is an e_mux
  assign p48_full_48 = ((read & !write) == 0)? full_47 :
    full_49;

  //control_reg_48, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_48 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_48 <= 0;
          else 
            full_48 <= p48_full_48;
    end


  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    stage_48;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    full_48;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_s1_arbitrator (
                                       // inputs:
                                        clk,
                                        cpu_data_master_address_to_slave,
                                        cpu_data_master_byteenable,
                                        cpu_data_master_debugaccess,
                                        cpu_data_master_latency_counter,
                                        cpu_data_master_read,
                                        cpu_data_master_write,
                                        cpu_data_master_writedata,
                                        cpu_instruction_master_address_to_slave,
                                        cpu_instruction_master_latency_counter,
                                        cpu_instruction_master_read,
                                        pipeline_bridge_s1_endofpacket,
                                        pipeline_bridge_s1_readdata,
                                        pipeline_bridge_s1_readdatavalid,
                                        pipeline_bridge_s1_waitrequest,
                                        reset_n,

                                       // outputs:
                                        cpu_data_master_granted_pipeline_bridge_s1,
                                        cpu_data_master_qualified_request_pipeline_bridge_s1,
                                        cpu_data_master_read_data_valid_pipeline_bridge_s1,
                                        cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
                                        cpu_data_master_requests_pipeline_bridge_s1,
                                        cpu_instruction_master_granted_pipeline_bridge_s1,
                                        cpu_instruction_master_qualified_request_pipeline_bridge_s1,
                                        cpu_instruction_master_read_data_valid_pipeline_bridge_s1,
                                        cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register,
                                        cpu_instruction_master_requests_pipeline_bridge_s1,
                                        d1_pipeline_bridge_s1_end_xfer,
                                        pipeline_bridge_s1_address,
                                        pipeline_bridge_s1_arbiterlock,
                                        pipeline_bridge_s1_arbiterlock2,
                                        pipeline_bridge_s1_burstcount,
                                        pipeline_bridge_s1_byteenable,
                                        pipeline_bridge_s1_chipselect,
                                        pipeline_bridge_s1_debugaccess,
                                        pipeline_bridge_s1_endofpacket_from_sa,
                                        pipeline_bridge_s1_nativeaddress,
                                        pipeline_bridge_s1_read,
                                        pipeline_bridge_s1_readdata_from_sa,
                                        pipeline_bridge_s1_reset_n,
                                        pipeline_bridge_s1_waitrequest_from_sa,
                                        pipeline_bridge_s1_write,
                                        pipeline_bridge_s1_writedata
                                     )
;

  output           cpu_data_master_granted_pipeline_bridge_s1;
  output           cpu_data_master_qualified_request_pipeline_bridge_s1;
  output           cpu_data_master_read_data_valid_pipeline_bridge_s1;
  output           cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register;
  output           cpu_data_master_requests_pipeline_bridge_s1;
  output           cpu_instruction_master_granted_pipeline_bridge_s1;
  output           cpu_instruction_master_qualified_request_pipeline_bridge_s1;
  output           cpu_instruction_master_read_data_valid_pipeline_bridge_s1;
  output           cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register;
  output           cpu_instruction_master_requests_pipeline_bridge_s1;
  output           d1_pipeline_bridge_s1_end_xfer;
  output  [ 24: 0] pipeline_bridge_s1_address;
  output           pipeline_bridge_s1_arbiterlock;
  output           pipeline_bridge_s1_arbiterlock2;
  output           pipeline_bridge_s1_burstcount;
  output  [  3: 0] pipeline_bridge_s1_byteenable;
  output           pipeline_bridge_s1_chipselect;
  output           pipeline_bridge_s1_debugaccess;
  output           pipeline_bridge_s1_endofpacket_from_sa;
  output  [ 24: 0] pipeline_bridge_s1_nativeaddress;
  output           pipeline_bridge_s1_read;
  output  [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  output           pipeline_bridge_s1_reset_n;
  output           pipeline_bridge_s1_waitrequest_from_sa;
  output           pipeline_bridge_s1_write;
  output  [ 31: 0] pipeline_bridge_s1_writedata;
  input            clk;
  input   [ 27: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 26: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            pipeline_bridge_s1_endofpacket;
  input   [ 31: 0] pipeline_bridge_s1_readdata;
  input            pipeline_bridge_s1_readdatavalid;
  input            pipeline_bridge_s1_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_pipeline_bridge_s1;
  wire             cpu_data_master_qualified_request_pipeline_bridge_s1;
  wire             cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1;
  wire             cpu_data_master_rdv_fifo_output_from_pipeline_bridge_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register;
  wire             cpu_data_master_requests_pipeline_bridge_s1;
  wire             cpu_data_master_saved_grant_pipeline_bridge_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_pipeline_bridge_s1;
  wire             cpu_instruction_master_qualified_request_pipeline_bridge_s1;
  wire             cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1;
  wire             cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register;
  wire             cpu_instruction_master_requests_pipeline_bridge_s1;
  wire             cpu_instruction_master_saved_grant_pipeline_bridge_s1;
  reg              d1_pipeline_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pipeline_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1;
  wire    [ 24: 0] pipeline_bridge_s1_address;
  wire             pipeline_bridge_s1_allgrants;
  wire             pipeline_bridge_s1_allow_new_arb_cycle;
  wire             pipeline_bridge_s1_any_bursting_master_saved_grant;
  wire             pipeline_bridge_s1_any_continuerequest;
  reg     [  1: 0] pipeline_bridge_s1_arb_addend;
  wire             pipeline_bridge_s1_arb_counter_enable;
  reg     [  3: 0] pipeline_bridge_s1_arb_share_counter;
  wire    [  3: 0] pipeline_bridge_s1_arb_share_counter_next_value;
  wire    [  3: 0] pipeline_bridge_s1_arb_share_set_values;
  wire    [  1: 0] pipeline_bridge_s1_arb_winner;
  wire             pipeline_bridge_s1_arbiterlock;
  wire             pipeline_bridge_s1_arbiterlock2;
  wire             pipeline_bridge_s1_arbitration_holdoff_internal;
  wire             pipeline_bridge_s1_beginbursttransfer_internal;
  wire             pipeline_bridge_s1_begins_xfer;
  wire             pipeline_bridge_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_s1_byteenable;
  wire             pipeline_bridge_s1_chipselect;
  wire    [  3: 0] pipeline_bridge_s1_chosen_master_double_vector;
  wire    [  1: 0] pipeline_bridge_s1_chosen_master_rot_left;
  wire             pipeline_bridge_s1_debugaccess;
  wire             pipeline_bridge_s1_end_xfer;
  wire             pipeline_bridge_s1_endofpacket_from_sa;
  wire             pipeline_bridge_s1_firsttransfer;
  wire    [  1: 0] pipeline_bridge_s1_grant_vector;
  wire             pipeline_bridge_s1_in_a_read_cycle;
  wire             pipeline_bridge_s1_in_a_write_cycle;
  wire    [  1: 0] pipeline_bridge_s1_master_qreq_vector;
  wire             pipeline_bridge_s1_move_on_to_next_transaction;
  wire    [ 24: 0] pipeline_bridge_s1_nativeaddress;
  wire             pipeline_bridge_s1_non_bursting_master_requests;
  wire             pipeline_bridge_s1_read;
  wire    [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  wire             pipeline_bridge_s1_readdatavalid_from_sa;
  reg              pipeline_bridge_s1_reg_firsttransfer;
  wire             pipeline_bridge_s1_reset_n;
  reg     [  1: 0] pipeline_bridge_s1_saved_chosen_master_vector;
  reg              pipeline_bridge_s1_slavearbiterlockenable;
  wire             pipeline_bridge_s1_slavearbiterlockenable2;
  wire             pipeline_bridge_s1_unreg_firsttransfer;
  wire             pipeline_bridge_s1_waitrequest_from_sa;
  wire             pipeline_bridge_s1_waits_for_read;
  wire             pipeline_bridge_s1_waits_for_write;
  wire             pipeline_bridge_s1_write;
  wire    [ 31: 0] pipeline_bridge_s1_writedata;
  wire    [ 27: 0] shifted_address_to_pipeline_bridge_s1_from_cpu_data_master;
  wire    [ 26: 0] shifted_address_to_pipeline_bridge_s1_from_cpu_instruction_master;
  wire             wait_for_pipeline_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pipeline_bridge_s1_end_xfer;
    end


  assign pipeline_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_pipeline_bridge_s1 | cpu_instruction_master_qualified_request_pipeline_bridge_s1));
  //assign pipeline_bridge_s1_readdatavalid_from_sa = pipeline_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_readdatavalid_from_sa = pipeline_bridge_s1_readdatavalid;

  //assign pipeline_bridge_s1_readdata_from_sa = pipeline_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_readdata_from_sa = pipeline_bridge_s1_readdata;

  assign cpu_data_master_requests_pipeline_bridge_s1 = ({cpu_data_master_address_to_slave[27] , 27'b0} == 28'h0) & (cpu_data_master_read | cpu_data_master_write);
  //assign pipeline_bridge_s1_waitrequest_from_sa = pipeline_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_waitrequest_from_sa = pipeline_bridge_s1_waitrequest;

  //pipeline_bridge_s1_arb_share_counter set values, which is an e_mux
  assign pipeline_bridge_s1_arb_share_set_values = (cpu_data_master_granted_pipeline_bridge_s1)? 8 :
    (cpu_instruction_master_granted_pipeline_bridge_s1)? 8 :
    (cpu_data_master_granted_pipeline_bridge_s1)? 8 :
    (cpu_instruction_master_granted_pipeline_bridge_s1)? 8 :
    (cpu_data_master_granted_pipeline_bridge_s1)? 8 :
    (cpu_instruction_master_granted_pipeline_bridge_s1)? 8 :
    1;

  //pipeline_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign pipeline_bridge_s1_non_bursting_master_requests = cpu_data_master_requests_pipeline_bridge_s1 |
    cpu_instruction_master_requests_pipeline_bridge_s1 |
    cpu_data_master_requests_pipeline_bridge_s1 |
    cpu_instruction_master_requests_pipeline_bridge_s1 |
    cpu_data_master_requests_pipeline_bridge_s1 |
    cpu_instruction_master_requests_pipeline_bridge_s1;

  //pipeline_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pipeline_bridge_s1_any_bursting_master_saved_grant = 0;

  //pipeline_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pipeline_bridge_s1_arb_share_counter_next_value = pipeline_bridge_s1_firsttransfer ? (pipeline_bridge_s1_arb_share_set_values - 1) : |pipeline_bridge_s1_arb_share_counter ? (pipeline_bridge_s1_arb_share_counter - 1) : 0;

  //pipeline_bridge_s1_allgrants all slave grants, which is an e_mux
  assign pipeline_bridge_s1_allgrants = (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector);

  //pipeline_bridge_s1_end_xfer assignment, which is an e_assign
  assign pipeline_bridge_s1_end_xfer = ~(pipeline_bridge_s1_waits_for_read | pipeline_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pipeline_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pipeline_bridge_s1 = pipeline_bridge_s1_end_xfer & (~pipeline_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pipeline_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pipeline_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pipeline_bridge_s1 & pipeline_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_pipeline_bridge_s1 & ~pipeline_bridge_s1_non_bursting_master_requests);

  //pipeline_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_arb_share_counter <= 0;
      else if (pipeline_bridge_s1_arb_counter_enable)
          pipeline_bridge_s1_arb_share_counter <= pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|pipeline_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pipeline_bridge_s1) | (end_xfer_arb_share_counter_term_pipeline_bridge_s1 & ~pipeline_bridge_s1_non_bursting_master_requests))
          pipeline_bridge_s1_slavearbiterlockenable <= |pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //cpu/data_master pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = pipeline_bridge_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //pipeline_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pipeline_bridge_s1_slavearbiterlockenable2 = |pipeline_bridge_s1_arb_share_counter_next_value;

  //cpu/data_master pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = pipeline_bridge_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = pipeline_bridge_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = pipeline_bridge_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 <= cpu_instruction_master_saved_grant_pipeline_bridge_s1 ? 1 : (pipeline_bridge_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_pipeline_bridge_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 & cpu_instruction_master_requests_pipeline_bridge_s1;

  //pipeline_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pipeline_bridge_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_pipeline_bridge_s1 = cpu_data_master_requests_pipeline_bridge_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter))) | cpu_instruction_master_arbiterlock);
  //unique name for pipeline_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign pipeline_bridge_s1_move_on_to_next_transaction = pipeline_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_pipeline_bridge_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1),
      .full                 (),
      .read                 (pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1;
  //local readdatavalid cpu_data_master_read_data_valid_pipeline_bridge_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_pipeline_bridge_s1 = (pipeline_bridge_s1_readdatavalid_from_sa & cpu_data_master_rdv_fifo_output_from_pipeline_bridge_s1) & ~ cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1;

  //pipeline_bridge_s1_writedata mux, which is an e_mux
  assign pipeline_bridge_s1_writedata = cpu_data_master_writedata;

  //assign pipeline_bridge_s1_endofpacket_from_sa = pipeline_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_endofpacket_from_sa = pipeline_bridge_s1_endofpacket;

  assign cpu_instruction_master_requests_pipeline_bridge_s1 = ((1) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 <= cpu_data_master_saved_grant_pipeline_bridge_s1 ? 1 : (pipeline_bridge_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_pipeline_bridge_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 & cpu_data_master_requests_pipeline_bridge_s1;

  assign cpu_instruction_master_qualified_request_pipeline_bridge_s1 = cpu_instruction_master_requests_pipeline_bridge_s1 & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter))) | cpu_data_master_arbiterlock);
  //rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_pipeline_bridge_s1),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1),
      .full                 (),
      .read                 (pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_s1_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register = ~cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1;
  //local readdatavalid cpu_instruction_master_read_data_valid_pipeline_bridge_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_pipeline_bridge_s1 = (pipeline_bridge_s1_readdatavalid_from_sa & cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_s1) & ~ cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1;

  //allow new arb cycle for pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_s1_master_qreq_vector[0] = cpu_instruction_master_qualified_request_pipeline_bridge_s1;

  //cpu/instruction_master grant pipeline_bridge/s1, which is an e_assign
  assign cpu_instruction_master_granted_pipeline_bridge_s1 = pipeline_bridge_s1_grant_vector[0];

  //cpu/instruction_master saved-grant pipeline_bridge/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_pipeline_bridge_s1 = pipeline_bridge_s1_arb_winner[0] && cpu_instruction_master_requests_pipeline_bridge_s1;

  //cpu/data_master assignment into master qualified-requests vector for pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_s1_master_qreq_vector[1] = cpu_data_master_qualified_request_pipeline_bridge_s1;

  //cpu/data_master grant pipeline_bridge/s1, which is an e_assign
  assign cpu_data_master_granted_pipeline_bridge_s1 = pipeline_bridge_s1_grant_vector[1];

  //cpu/data_master saved-grant pipeline_bridge/s1, which is an e_assign
  assign cpu_data_master_saved_grant_pipeline_bridge_s1 = pipeline_bridge_s1_arb_winner[1] && cpu_data_master_requests_pipeline_bridge_s1;

  //pipeline_bridge/s1 chosen-master double-vector, which is an e_assign
  assign pipeline_bridge_s1_chosen_master_double_vector = {pipeline_bridge_s1_master_qreq_vector, pipeline_bridge_s1_master_qreq_vector} & ({~pipeline_bridge_s1_master_qreq_vector, ~pipeline_bridge_s1_master_qreq_vector} + pipeline_bridge_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pipeline_bridge_s1_arb_winner = (pipeline_bridge_s1_allow_new_arb_cycle & | pipeline_bridge_s1_grant_vector) ? pipeline_bridge_s1_grant_vector : pipeline_bridge_s1_saved_chosen_master_vector;

  //saved pipeline_bridge_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_saved_chosen_master_vector <= 0;
      else if (pipeline_bridge_s1_allow_new_arb_cycle)
          pipeline_bridge_s1_saved_chosen_master_vector <= |pipeline_bridge_s1_grant_vector ? pipeline_bridge_s1_grant_vector : pipeline_bridge_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pipeline_bridge_s1_grant_vector = {(pipeline_bridge_s1_chosen_master_double_vector[1] | pipeline_bridge_s1_chosen_master_double_vector[3]),
    (pipeline_bridge_s1_chosen_master_double_vector[0] | pipeline_bridge_s1_chosen_master_double_vector[2])};

  //pipeline_bridge/s1 chosen master rotated left, which is an e_assign
  assign pipeline_bridge_s1_chosen_master_rot_left = (pipeline_bridge_s1_arb_winner << 1) ? (pipeline_bridge_s1_arb_winner << 1) : 1;

  //pipeline_bridge/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_arb_addend <= 1;
      else if (|pipeline_bridge_s1_grant_vector)
          pipeline_bridge_s1_arb_addend <= pipeline_bridge_s1_end_xfer? pipeline_bridge_s1_chosen_master_rot_left : pipeline_bridge_s1_grant_vector;
    end


  //pipeline_bridge_s1_reset_n assignment, which is an e_assign
  assign pipeline_bridge_s1_reset_n = reset_n;

  assign pipeline_bridge_s1_chipselect = cpu_data_master_granted_pipeline_bridge_s1 | cpu_instruction_master_granted_pipeline_bridge_s1;
  //pipeline_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_s1_firsttransfer = pipeline_bridge_s1_begins_xfer ? pipeline_bridge_s1_unreg_firsttransfer : pipeline_bridge_s1_reg_firsttransfer;

  //pipeline_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_s1_unreg_firsttransfer = ~(pipeline_bridge_s1_slavearbiterlockenable & pipeline_bridge_s1_any_continuerequest);

  //pipeline_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (pipeline_bridge_s1_begins_xfer)
          pipeline_bridge_s1_reg_firsttransfer <= pipeline_bridge_s1_unreg_firsttransfer;
    end


  //pipeline_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pipeline_bridge_s1_beginbursttransfer_internal = pipeline_bridge_s1_begins_xfer;

  //pipeline_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pipeline_bridge_s1_arbitration_holdoff_internal = pipeline_bridge_s1_begins_xfer & pipeline_bridge_s1_firsttransfer;

  //pipeline_bridge_s1_read assignment, which is an e_mux
  assign pipeline_bridge_s1_read = (cpu_data_master_granted_pipeline_bridge_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pipeline_bridge_s1 & cpu_instruction_master_read);

  //pipeline_bridge_s1_write assignment, which is an e_mux
  assign pipeline_bridge_s1_write = cpu_data_master_granted_pipeline_bridge_s1 & cpu_data_master_write;

  assign shifted_address_to_pipeline_bridge_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //pipeline_bridge_s1_address mux, which is an e_mux
  assign pipeline_bridge_s1_address = (cpu_data_master_granted_pipeline_bridge_s1)? (shifted_address_to_pipeline_bridge_s1_from_cpu_data_master >> 2) :
    (shifted_address_to_pipeline_bridge_s1_from_cpu_instruction_master >> 2);

  assign shifted_address_to_pipeline_bridge_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //slaveid pipeline_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pipeline_bridge_s1_nativeaddress = (cpu_data_master_granted_pipeline_bridge_s1)? (cpu_data_master_address_to_slave >> 2) :
    (cpu_instruction_master_address_to_slave >> 2);

  //d1_pipeline_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pipeline_bridge_s1_end_xfer <= 1;
      else 
        d1_pipeline_bridge_s1_end_xfer <= pipeline_bridge_s1_end_xfer;
    end


  //pipeline_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign pipeline_bridge_s1_waits_for_read = pipeline_bridge_s1_in_a_read_cycle & pipeline_bridge_s1_waitrequest_from_sa;

  //pipeline_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign pipeline_bridge_s1_in_a_read_cycle = (cpu_data_master_granted_pipeline_bridge_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pipeline_bridge_s1 & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pipeline_bridge_s1_in_a_read_cycle;

  //pipeline_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign pipeline_bridge_s1_waits_for_write = pipeline_bridge_s1_in_a_write_cycle & pipeline_bridge_s1_waitrequest_from_sa;

  //pipeline_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign pipeline_bridge_s1_in_a_write_cycle = cpu_data_master_granted_pipeline_bridge_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pipeline_bridge_s1_in_a_write_cycle;

  assign wait_for_pipeline_bridge_s1_counter = 0;
  //pipeline_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign pipeline_bridge_s1_byteenable = (cpu_data_master_granted_pipeline_bridge_s1)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pipeline_bridge_s1_burstcount = 1;

  //pipeline_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pipeline_bridge_s1_arbiterlock = (cpu_data_master_arbiterlock)? cpu_data_master_arbiterlock :
    cpu_instruction_master_arbiterlock;

  //pipeline_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pipeline_bridge_s1_arbiterlock2 = (cpu_data_master_arbiterlock2)? cpu_data_master_arbiterlock2 :
    cpu_instruction_master_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pipeline_bridge_s1_debugaccess = (cpu_data_master_granted_pipeline_bridge_s1)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_pipeline_bridge_s1 + cpu_instruction_master_granted_pipeline_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_pipeline_bridge_s1 + cpu_instruction_master_saved_grant_pipeline_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_module (
                                                                                      // inputs:
                                                                                       clear_fifo,
                                                                                       clk,
                                                                                       data_in,
                                                                                       read,
                                                                                       reset_n,
                                                                                       sync_reset,
                                                                                       write,

                                                                                      // outputs:
                                                                                       data_out,
                                                                                       empty,
                                                                                       fifo_contains_ones_n,
                                                                                       full
                                                                                    )
;

  output  [  2: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  2: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  2: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  2: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  2: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  2: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  2: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  2: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  2: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  2: 0] p6_stage_6;
  reg     [  2: 0] stage_0;
  reg     [  2: 0] stage_1;
  reg     [  2: 0] stage_2;
  reg     [  2: 0] stage_3;
  reg     [  2: 0] stage_4;
  reg     [  2: 0] stage_5;
  reg     [  2: 0] stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_m1_arbitrator (
                                       // inputs:
                                        clk,
                                        clock_crossing_bridge_s1_endofpacket_from_sa,
                                        clock_crossing_bridge_s1_readdata_from_sa,
                                        clock_crossing_bridge_s1_waitrequest_from_sa,
                                        colour_lookup_table_s1_readdata_from_sa,
                                        cpu_jtag_debug_module_readdata_from_sa,
                                        d1_clock_crossing_bridge_s1_end_xfer,
                                        d1_colour_lookup_table_s1_end_xfer,
                                        d1_cpu_jtag_debug_module_end_xfer,
                                        d1_descriptor_memory_s1_end_xfer,
                                        d1_flash_ssram_pipeline_bridge_s1_end_xfer,
                                        d1_frame_buffer_pipeline_bridge_s1_end_xfer,
                                        d1_lcd_sgdma_csr_end_xfer,
                                        descriptor_memory_s1_readdata_from_sa,
                                        flash_ssram_pipeline_bridge_s1_endofpacket_from_sa,
                                        flash_ssram_pipeline_bridge_s1_readdata_from_sa,
                                        flash_ssram_pipeline_bridge_s1_waitrequest_from_sa,
                                        frame_buffer_pipeline_bridge_s1_endofpacket_from_sa,
                                        frame_buffer_pipeline_bridge_s1_readdata_from_sa,
                                        frame_buffer_pipeline_bridge_s1_waitrequest_from_sa,
                                        lcd_sgdma_csr_readdata_from_sa,
                                        pipeline_bridge_m1_address,
                                        pipeline_bridge_m1_burstcount,
                                        pipeline_bridge_m1_byteenable,
                                        pipeline_bridge_m1_chipselect,
                                        pipeline_bridge_m1_granted_clock_crossing_bridge_s1,
                                        pipeline_bridge_m1_granted_colour_lookup_table_s1,
                                        pipeline_bridge_m1_granted_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_granted_descriptor_memory_s1,
                                        pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1,
                                        pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1,
                                        pipeline_bridge_m1_granted_lcd_sgdma_csr,
                                        pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1,
                                        pipeline_bridge_m1_qualified_request_colour_lookup_table_s1,
                                        pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_qualified_request_descriptor_memory_s1,
                                        pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1,
                                        pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1,
                                        pipeline_bridge_m1_qualified_request_lcd_sgdma_csr,
                                        pipeline_bridge_m1_read,
                                        pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1,
                                        pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register,
                                        pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1,
                                        pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_read_data_valid_descriptor_memory_s1,
                                        pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1,
                                        pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
                                        pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1,
                                        pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register,
                                        pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr,
                                        pipeline_bridge_m1_requests_clock_crossing_bridge_s1,
                                        pipeline_bridge_m1_requests_colour_lookup_table_s1,
                                        pipeline_bridge_m1_requests_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_requests_descriptor_memory_s1,
                                        pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1,
                                        pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1,
                                        pipeline_bridge_m1_requests_lcd_sgdma_csr,
                                        pipeline_bridge_m1_write,
                                        pipeline_bridge_m1_writedata,
                                        reset_n,

                                       // outputs:
                                        pipeline_bridge_m1_address_to_slave,
                                        pipeline_bridge_m1_endofpacket,
                                        pipeline_bridge_m1_latency_counter,
                                        pipeline_bridge_m1_readdata,
                                        pipeline_bridge_m1_readdatavalid,
                                        pipeline_bridge_m1_waitrequest
                                     )
;

  output  [ 26: 0] pipeline_bridge_m1_address_to_slave;
  output           pipeline_bridge_m1_endofpacket;
  output           pipeline_bridge_m1_latency_counter;
  output  [ 31: 0] pipeline_bridge_m1_readdata;
  output           pipeline_bridge_m1_readdatavalid;
  output           pipeline_bridge_m1_waitrequest;
  input            clk;
  input            clock_crossing_bridge_s1_endofpacket_from_sa;
  input   [ 31: 0] clock_crossing_bridge_s1_readdata_from_sa;
  input            clock_crossing_bridge_s1_waitrequest_from_sa;
  input   [ 31: 0] colour_lookup_table_s1_readdata_from_sa;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_clock_crossing_bridge_s1_end_xfer;
  input            d1_colour_lookup_table_s1_end_xfer;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_descriptor_memory_s1_end_xfer;
  input            d1_flash_ssram_pipeline_bridge_s1_end_xfer;
  input            d1_frame_buffer_pipeline_bridge_s1_end_xfer;
  input            d1_lcd_sgdma_csr_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            flash_ssram_pipeline_bridge_s1_endofpacket_from_sa;
  input   [255: 0] flash_ssram_pipeline_bridge_s1_readdata_from_sa;
  input            flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
  input            frame_buffer_pipeline_bridge_s1_endofpacket_from_sa;
  input   [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata_from_sa;
  input            frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;
  input   [ 31: 0] lcd_sgdma_csr_readdata_from_sa;
  input   [ 26: 0] pipeline_bridge_m1_address;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_granted_clock_crossing_bridge_s1;
  input            pipeline_bridge_m1_granted_colour_lookup_table_s1;
  input            pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_granted_descriptor_memory_s1;
  input            pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1;
  input            pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1;
  input            pipeline_bridge_m1_granted_lcd_sgdma_csr;
  input            pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1;
  input            pipeline_bridge_m1_qualified_request_colour_lookup_table_s1;
  input            pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_qualified_request_descriptor_memory_s1;
  input            pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1;
  input            pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1;
  input            pipeline_bridge_m1_qualified_request_lcd_sgdma_csr;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1;
  input            pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1;
  input            pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_read_data_valid_descriptor_memory_s1;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1;
  input            pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1;
  input            pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  input            pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr;
  input            pipeline_bridge_m1_requests_clock_crossing_bridge_s1;
  input            pipeline_bridge_m1_requests_colour_lookup_table_s1;
  input            pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_requests_descriptor_memory_s1;
  input            pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;
  input            pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1;
  input            pipeline_bridge_m1_requests_lcd_sgdma_csr;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             empty_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo;
  wire    [ 31: 0] flash_ssram_pipeline_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs;
  wire             full_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo;
  wire             latency_load_value;
  wire             p1_pipeline_bridge_m1_latency_counter;
  reg     [ 26: 0] pipeline_bridge_m1_address_last_time;
  wire    [ 26: 0] pipeline_bridge_m1_address_to_slave;
  reg              pipeline_bridge_m1_burstcount_last_time;
  reg     [  3: 0] pipeline_bridge_m1_byteenable_last_time;
  reg              pipeline_bridge_m1_chipselect_last_time;
  wire             pipeline_bridge_m1_endofpacket;
  wire             pipeline_bridge_m1_is_granted_some_slave;
  reg              pipeline_bridge_m1_latency_counter;
  reg              pipeline_bridge_m1_read_but_no_slave_selected;
  reg              pipeline_bridge_m1_read_last_time;
  wire    [ 31: 0] pipeline_bridge_m1_readdata;
  wire             pipeline_bridge_m1_readdatavalid;
  wire             pipeline_bridge_m1_run;
  wire             pipeline_bridge_m1_waitrequest;
  reg              pipeline_bridge_m1_write_last_time;
  reg     [ 31: 0] pipeline_bridge_m1_writedata_last_time;
  wire             pre_flush_pipeline_bridge_m1_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             read_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo;
  wire    [  2: 0] selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output;
  wire    [  2: 0] selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1;
  wire             write_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1 | ~pipeline_bridge_m1_requests_clock_crossing_bridge_s1) & ((~pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1 | ~pipeline_bridge_m1_chipselect | (1 & ~clock_crossing_bridge_s1_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1 | ~pipeline_bridge_m1_chipselect | (1 & ~clock_crossing_bridge_s1_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_colour_lookup_table_s1 | ~pipeline_bridge_m1_requests_colour_lookup_table_s1) & ((~pipeline_bridge_m1_qualified_request_colour_lookup_table_s1 | ~pipeline_bridge_m1_chipselect | (1 & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_colour_lookup_table_s1 | ~pipeline_bridge_m1_chipselect | (1 & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module | ~pipeline_bridge_m1_requests_cpu_jtag_debug_module) & ((~pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module | ~(pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) | (1 & ~d1_cpu_jtag_debug_module_end_xfer & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))) & ((~pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module | ~(pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect) | (1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect)))) & 1 & (pipeline_bridge_m1_qualified_request_descriptor_memory_s1 | ~pipeline_bridge_m1_requests_descriptor_memory_s1) & ((~pipeline_bridge_m1_qualified_request_descriptor_memory_s1 | ~pipeline_bridge_m1_chipselect | (1 & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_descriptor_memory_s1 | ~pipeline_bridge_m1_chipselect | (1 & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1 | ~pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1) & ((~pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1 | ~pipeline_bridge_m1_chipselect | (1 & ~flash_ssram_pipeline_bridge_s1_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1 | ~pipeline_bridge_m1_chipselect | (1 & ~flash_ssram_pipeline_bridge_s1_waitrequest_from_sa & pipeline_bridge_m1_chipselect)));

  //cascaded wait assignment, which is an e_assign
  assign pipeline_bridge_m1_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1 | ~pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1) & (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 | ~pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1) & ((~pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1 | ~pipeline_bridge_m1_chipselect | (1 & ~frame_buffer_pipeline_bridge_s1_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1 | ~pipeline_bridge_m1_chipselect | (1 & ~frame_buffer_pipeline_bridge_s1_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_lcd_sgdma_csr | ~pipeline_bridge_m1_requests_lcd_sgdma_csr) & ((~pipeline_bridge_m1_qualified_request_lcd_sgdma_csr | ~(pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) | (1 & ~d1_lcd_sgdma_csr_end_xfer & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))) & ((~pipeline_bridge_m1_qualified_request_lcd_sgdma_csr | ~(pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect) | (1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect))));

  //optimize select-logic by passing only those address bits which matter.
  assign pipeline_bridge_m1_address_to_slave = pipeline_bridge_m1_address[26 : 0];

  //pipeline_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_but_no_slave_selected <= 0;
      else 
        pipeline_bridge_m1_read_but_no_slave_selected <= (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & pipeline_bridge_m1_run & ~pipeline_bridge_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pipeline_bridge_m1_is_granted_some_slave = pipeline_bridge_m1_granted_clock_crossing_bridge_s1 |
    pipeline_bridge_m1_granted_colour_lookup_table_s1 |
    pipeline_bridge_m1_granted_cpu_jtag_debug_module |
    pipeline_bridge_m1_granted_descriptor_memory_s1 |
    pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1 |
    pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1 |
    pipeline_bridge_m1_granted_lcd_sgdma_csr;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pipeline_bridge_m1_readdatavalid = pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1 |
    pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1 |
    pipeline_bridge_m1_read_data_valid_descriptor_memory_s1 |
    pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1 |
    pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pipeline_bridge_m1_readdatavalid = pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr;

  //pipeline_bridge/m1 readdata mux, which is an e_mux
  assign pipeline_bridge_m1_readdata = ({32 {~pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1}} | clock_crossing_bridge_s1_readdata_from_sa) &
    ({32 {~pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1}} | colour_lookup_table_s1_readdata_from_sa) &
    ({32 {~((pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~pipeline_bridge_m1_read_data_valid_descriptor_memory_s1}} | descriptor_memory_s1_readdata_from_sa) &
    ({32 {~pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1}} | flash_ssram_pipeline_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs) &
    ({32 {~pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1}} | frame_buffer_pipeline_bridge_s1_readdata_from_sa) &
    ({32 {~((pipeline_bridge_m1_qualified_request_lcd_sgdma_csr & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | lcd_sgdma_csr_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign pipeline_bridge_m1_waitrequest = ~pipeline_bridge_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_latency_counter <= 0;
      else 
        pipeline_bridge_m1_latency_counter <= p1_pipeline_bridge_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pipeline_bridge_m1_latency_counter = ((pipeline_bridge_m1_run & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))? latency_load_value :
    (pipeline_bridge_m1_latency_counter)? pipeline_bridge_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {pipeline_bridge_m1_requests_colour_lookup_table_s1}} & 1) |
    ({1 {pipeline_bridge_m1_requests_descriptor_memory_s1}} & 1);

  //mux pipeline_bridge_m1_endofpacket, which is an e_mux
  assign pipeline_bridge_m1_endofpacket = (pipeline_bridge_m1_requests_clock_crossing_bridge_s1)? clock_crossing_bridge_s1_endofpacket_from_sa :
    (pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1)? flash_ssram_pipeline_bridge_s1_endofpacket_from_sa :
    frame_buffer_pipeline_bridge_s1_endofpacket_from_sa;

  //Negative Dynamic Bus-sizing mux.
  //this mux selects the correct eighth of the 
  //wide data coming from the slave flash_ssram_pipeline_bridge/s1 
  assign flash_ssram_pipeline_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs = ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 0))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[31 : 0] :
    ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 1))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[63 : 32] :
    ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 2))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[95 : 64] :
    ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 3))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[127 : 96] :
    ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 4))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[159 : 128] :
    ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 5))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[191 : 160] :
    ((selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 == 6))? flash_ssram_pipeline_bridge_s1_readdata_from_sa[223 : 192] :
    flash_ssram_pipeline_bridge_s1_readdata_from_sa[255 : 224];

  //read_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo fifo read, which is an e_mux
  assign read_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo = pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1;

  //write_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo fifo write, which is an e_mux
  assign write_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo = (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & pipeline_bridge_m1_run & pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;

  assign selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output_flash_ssram_pipeline_bridge_s1 = selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output;
  //selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_module selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (pipeline_bridge_m1_address_to_slave[4 : 2]),
      .data_out             (selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo_output),
      .empty                (empty_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo),
      .fifo_contains_ones_n (),
      .full                 (full_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo),
      .read                 (read_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (write_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo)
    );


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_address_last_time <= 0;
      else 
        pipeline_bridge_m1_address_last_time <= pipeline_bridge_m1_address;
    end


  //pipeline_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pipeline_bridge_m1_waitrequest & pipeline_bridge_m1_chipselect;
    end


  //pipeline_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_address != pipeline_bridge_m1_address_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_chipselect_last_time <= 0;
      else 
        pipeline_bridge_m1_chipselect_last_time <= pipeline_bridge_m1_chipselect;
    end


  //pipeline_bridge_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_chipselect != pipeline_bridge_m1_chipselect_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_burstcount_last_time <= 0;
      else 
        pipeline_bridge_m1_burstcount_last_time <= pipeline_bridge_m1_burstcount;
    end


  //pipeline_bridge_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_burstcount != pipeline_bridge_m1_burstcount_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_byteenable_last_time <= 0;
      else 
        pipeline_bridge_m1_byteenable_last_time <= pipeline_bridge_m1_byteenable;
    end


  //pipeline_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_byteenable != pipeline_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_last_time <= 0;
      else 
        pipeline_bridge_m1_read_last_time <= pipeline_bridge_m1_read;
    end


  //pipeline_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_read != pipeline_bridge_m1_read_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_write_last_time <= 0;
      else 
        pipeline_bridge_m1_write_last_time <= pipeline_bridge_m1_write;
    end


  //pipeline_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_write != pipeline_bridge_m1_write_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_writedata_last_time <= 0;
      else 
        pipeline_bridge_m1_writedata_last_time <= pipeline_bridge_m1_writedata;
    end


  //pipeline_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_writedata != pipeline_bridge_m1_writedata_last_time) & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect))
        begin
          $write("%0d ns: pipeline_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end


  //selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo read when empty, which is an e_process
  always @(posedge clk)
    begin
      if (empty_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo & read_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo)
        begin
          $write("%0d ns: pipeline_bridge/m1 negative rdv fifo selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo: read AND empty.\n", $time);
          $stop;
        end
    end


  //selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo write when full, which is an e_process
  always @(posedge clk)
    begin
      if (full_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo & write_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo & ~read_selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo)
        begin
          $write("%0d ns: pipeline_bridge/m1 negative rdv fifo selecto_nrdv_pipeline_bridge_m1_3_flash_ssram_pipeline_bridge_s1_fifo: write AND full.\n", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module push_buttons_s1_arbitrator (
                                    // inputs:
                                     clk,
                                     clock_crossing_bridge_m1_address_to_slave,
                                     clock_crossing_bridge_m1_latency_counter,
                                     clock_crossing_bridge_m1_nativeaddress,
                                     clock_crossing_bridge_m1_read,
                                     clock_crossing_bridge_m1_write,
                                     clock_crossing_bridge_m1_writedata,
                                     push_buttons_s1_irq,
                                     push_buttons_s1_readdata,
                                     reset_n,

                                    // outputs:
                                     clock_crossing_bridge_m1_granted_push_buttons_s1,
                                     clock_crossing_bridge_m1_qualified_request_push_buttons_s1,
                                     clock_crossing_bridge_m1_read_data_valid_push_buttons_s1,
                                     clock_crossing_bridge_m1_requests_push_buttons_s1,
                                     d1_push_buttons_s1_end_xfer,
                                     push_buttons_s1_address,
                                     push_buttons_s1_chipselect,
                                     push_buttons_s1_irq_from_sa,
                                     push_buttons_s1_readdata_from_sa,
                                     push_buttons_s1_reset_n,
                                     push_buttons_s1_write_n,
                                     push_buttons_s1_writedata
                                  )
;

  output           clock_crossing_bridge_m1_granted_push_buttons_s1;
  output           clock_crossing_bridge_m1_qualified_request_push_buttons_s1;
  output           clock_crossing_bridge_m1_read_data_valid_push_buttons_s1;
  output           clock_crossing_bridge_m1_requests_push_buttons_s1;
  output           d1_push_buttons_s1_end_xfer;
  output  [  1: 0] push_buttons_s1_address;
  output           push_buttons_s1_chipselect;
  output           push_buttons_s1_irq_from_sa;
  output  [ 31: 0] push_buttons_s1_readdata_from_sa;
  output           push_buttons_s1_reset_n;
  output           push_buttons_s1_write_n;
  output  [ 31: 0] push_buttons_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input            push_buttons_s1_irq;
  input   [ 31: 0] push_buttons_s1_readdata;
  input            reset_n;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_push_buttons_s1;
  wire             clock_crossing_bridge_m1_qualified_request_push_buttons_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_push_buttons_s1;
  wire             clock_crossing_bridge_m1_requests_push_buttons_s1;
  wire             clock_crossing_bridge_m1_saved_grant_push_buttons_s1;
  reg              d1_push_buttons_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_push_buttons_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] push_buttons_s1_address;
  wire             push_buttons_s1_allgrants;
  wire             push_buttons_s1_allow_new_arb_cycle;
  wire             push_buttons_s1_any_bursting_master_saved_grant;
  wire             push_buttons_s1_any_continuerequest;
  wire             push_buttons_s1_arb_counter_enable;
  reg              push_buttons_s1_arb_share_counter;
  wire             push_buttons_s1_arb_share_counter_next_value;
  wire             push_buttons_s1_arb_share_set_values;
  wire             push_buttons_s1_beginbursttransfer_internal;
  wire             push_buttons_s1_begins_xfer;
  wire             push_buttons_s1_chipselect;
  wire             push_buttons_s1_end_xfer;
  wire             push_buttons_s1_firsttransfer;
  wire             push_buttons_s1_grant_vector;
  wire             push_buttons_s1_in_a_read_cycle;
  wire             push_buttons_s1_in_a_write_cycle;
  wire             push_buttons_s1_irq_from_sa;
  wire             push_buttons_s1_master_qreq_vector;
  wire             push_buttons_s1_non_bursting_master_requests;
  wire    [ 31: 0] push_buttons_s1_readdata_from_sa;
  reg              push_buttons_s1_reg_firsttransfer;
  wire             push_buttons_s1_reset_n;
  reg              push_buttons_s1_slavearbiterlockenable;
  wire             push_buttons_s1_slavearbiterlockenable2;
  wire             push_buttons_s1_unreg_firsttransfer;
  wire             push_buttons_s1_waits_for_read;
  wire             push_buttons_s1_waits_for_write;
  wire             push_buttons_s1_write_n;
  wire    [ 31: 0] push_buttons_s1_writedata;
  wire             wait_for_push_buttons_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~push_buttons_s1_end_xfer;
    end


  assign push_buttons_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_push_buttons_s1));
  //assign push_buttons_s1_readdata_from_sa = push_buttons_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign push_buttons_s1_readdata_from_sa = push_buttons_s1_readdata;

  assign clock_crossing_bridge_m1_requests_push_buttons_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h200) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //push_buttons_s1_arb_share_counter set values, which is an e_mux
  assign push_buttons_s1_arb_share_set_values = 1;

  //push_buttons_s1_non_bursting_master_requests mux, which is an e_mux
  assign push_buttons_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_push_buttons_s1;

  //push_buttons_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign push_buttons_s1_any_bursting_master_saved_grant = 0;

  //push_buttons_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign push_buttons_s1_arb_share_counter_next_value = push_buttons_s1_firsttransfer ? (push_buttons_s1_arb_share_set_values - 1) : |push_buttons_s1_arb_share_counter ? (push_buttons_s1_arb_share_counter - 1) : 0;

  //push_buttons_s1_allgrants all slave grants, which is an e_mux
  assign push_buttons_s1_allgrants = |push_buttons_s1_grant_vector;

  //push_buttons_s1_end_xfer assignment, which is an e_assign
  assign push_buttons_s1_end_xfer = ~(push_buttons_s1_waits_for_read | push_buttons_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_push_buttons_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_push_buttons_s1 = push_buttons_s1_end_xfer & (~push_buttons_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //push_buttons_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign push_buttons_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_push_buttons_s1 & push_buttons_s1_allgrants) | (end_xfer_arb_share_counter_term_push_buttons_s1 & ~push_buttons_s1_non_bursting_master_requests);

  //push_buttons_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          push_buttons_s1_arb_share_counter <= 0;
      else if (push_buttons_s1_arb_counter_enable)
          push_buttons_s1_arb_share_counter <= push_buttons_s1_arb_share_counter_next_value;
    end


  //push_buttons_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          push_buttons_s1_slavearbiterlockenable <= 0;
      else if ((|push_buttons_s1_master_qreq_vector & end_xfer_arb_share_counter_term_push_buttons_s1) | (end_xfer_arb_share_counter_term_push_buttons_s1 & ~push_buttons_s1_non_bursting_master_requests))
          push_buttons_s1_slavearbiterlockenable <= |push_buttons_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 push_buttons/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = push_buttons_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //push_buttons_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign push_buttons_s1_slavearbiterlockenable2 = |push_buttons_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 push_buttons/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = push_buttons_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //push_buttons_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign push_buttons_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_push_buttons_s1 = clock_crossing_bridge_m1_requests_push_buttons_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_push_buttons_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_push_buttons_s1 = clock_crossing_bridge_m1_granted_push_buttons_s1 & clock_crossing_bridge_m1_read & ~push_buttons_s1_waits_for_read;

  //push_buttons_s1_writedata mux, which is an e_mux
  assign push_buttons_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_push_buttons_s1 = clock_crossing_bridge_m1_qualified_request_push_buttons_s1;

  //clock_crossing_bridge/m1 saved-grant push_buttons/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_push_buttons_s1 = clock_crossing_bridge_m1_requests_push_buttons_s1;

  //allow new arb cycle for push_buttons/s1, which is an e_assign
  assign push_buttons_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign push_buttons_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign push_buttons_s1_master_qreq_vector = 1;

  //push_buttons_s1_reset_n assignment, which is an e_assign
  assign push_buttons_s1_reset_n = reset_n;

  assign push_buttons_s1_chipselect = clock_crossing_bridge_m1_granted_push_buttons_s1;
  //push_buttons_s1_firsttransfer first transaction, which is an e_assign
  assign push_buttons_s1_firsttransfer = push_buttons_s1_begins_xfer ? push_buttons_s1_unreg_firsttransfer : push_buttons_s1_reg_firsttransfer;

  //push_buttons_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign push_buttons_s1_unreg_firsttransfer = ~(push_buttons_s1_slavearbiterlockenable & push_buttons_s1_any_continuerequest);

  //push_buttons_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          push_buttons_s1_reg_firsttransfer <= 1'b1;
      else if (push_buttons_s1_begins_xfer)
          push_buttons_s1_reg_firsttransfer <= push_buttons_s1_unreg_firsttransfer;
    end


  //push_buttons_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign push_buttons_s1_beginbursttransfer_internal = push_buttons_s1_begins_xfer;

  //~push_buttons_s1_write_n assignment, which is an e_mux
  assign push_buttons_s1_write_n = ~(clock_crossing_bridge_m1_granted_push_buttons_s1 & clock_crossing_bridge_m1_write);

  //push_buttons_s1_address mux, which is an e_mux
  assign push_buttons_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_push_buttons_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_push_buttons_s1_end_xfer <= 1;
      else 
        d1_push_buttons_s1_end_xfer <= push_buttons_s1_end_xfer;
    end


  //push_buttons_s1_waits_for_read in a cycle, which is an e_mux
  assign push_buttons_s1_waits_for_read = push_buttons_s1_in_a_read_cycle & push_buttons_s1_begins_xfer;

  //push_buttons_s1_in_a_read_cycle assignment, which is an e_assign
  assign push_buttons_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_push_buttons_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = push_buttons_s1_in_a_read_cycle;

  //push_buttons_s1_waits_for_write in a cycle, which is an e_mux
  assign push_buttons_s1_waits_for_write = push_buttons_s1_in_a_write_cycle & 0;

  //push_buttons_s1_in_a_write_cycle assignment, which is an e_assign
  assign push_buttons_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_push_buttons_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = push_buttons_s1_in_a_write_cycle;

  assign wait_for_push_buttons_s1_counter = 0;
  //assign push_buttons_s1_irq_from_sa = push_buttons_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign push_buttons_s1_irq_from_sa = push_buttons_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //push_buttons/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         clock_crossing_bridge_m1_address_to_slave,
                                         clock_crossing_bridge_m1_latency_counter,
                                         clock_crossing_bridge_m1_nativeaddress,
                                         clock_crossing_bridge_m1_read,
                                         clock_crossing_bridge_m1_write,
                                         reset_n,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         clock_crossing_bridge_m1_granted_sysid_control_slave,
                                         clock_crossing_bridge_m1_qualified_request_sysid_control_slave,
                                         clock_crossing_bridge_m1_read_data_valid_sysid_control_slave,
                                         clock_crossing_bridge_m1_requests_sysid_control_slave,
                                         d1_sysid_control_slave_end_xfer,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa,
                                         sysid_control_slave_reset_n
                                      )
;

  output           clock_crossing_bridge_m1_granted_sysid_control_slave;
  output           clock_crossing_bridge_m1_qualified_request_sysid_control_slave;
  output           clock_crossing_bridge_m1_read_data_valid_sysid_control_slave;
  output           clock_crossing_bridge_m1_requests_sysid_control_slave;
  output           d1_sysid_control_slave_end_xfer;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  output           sysid_control_slave_reset_n;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_sysid_control_slave;
  wire             clock_crossing_bridge_m1_qualified_request_sysid_control_slave;
  wire             clock_crossing_bridge_m1_read_data_valid_sysid_control_slave;
  wire             clock_crossing_bridge_m1_requests_sysid_control_slave;
  wire             clock_crossing_bridge_m1_saved_grant_sysid_control_slave;
  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg              sysid_control_slave_arb_share_counter;
  wire             sysid_control_slave_arb_share_counter_next_value;
  wire             sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  wire             sysid_control_slave_reset_n;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign clock_crossing_bridge_m1_requests_sysid_control_slave = (({clock_crossing_bridge_m1_address_to_slave[10 : 3] , 3'b0} == 11'h5c0) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write)) & clock_crossing_bridge_m1_read;
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = clock_crossing_bridge_m1_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 sysid/control_slave arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = sysid_control_slave_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 sysid/control_slave arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_sysid_control_slave = clock_crossing_bridge_m1_requests_sysid_control_slave & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_sysid_control_slave, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_sysid_control_slave = clock_crossing_bridge_m1_granted_sysid_control_slave & clock_crossing_bridge_m1_read & ~sysid_control_slave_waits_for_read;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_sysid_control_slave = clock_crossing_bridge_m1_qualified_request_sysid_control_slave;

  //clock_crossing_bridge/m1 saved-grant sysid/control_slave, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_sysid_control_slave = clock_crossing_bridge_m1_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_reset_n assignment, which is an e_assign
  assign sysid_control_slave_reset_n = reset_n;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = clock_crossing_bridge_m1_granted_sysid_control_slave & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = clock_crossing_bridge_m1_granted_sysid_control_slave & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_tick_s1_arbitrator (
                                   // inputs:
                                    clk,
                                    clock_crossing_bridge_m1_address_to_slave,
                                    clock_crossing_bridge_m1_latency_counter,
                                    clock_crossing_bridge_m1_nativeaddress,
                                    clock_crossing_bridge_m1_read,
                                    clock_crossing_bridge_m1_write,
                                    clock_crossing_bridge_m1_writedata,
                                    reset_n,
                                    system_tick_s1_irq,
                                    system_tick_s1_readdata,

                                   // outputs:
                                    clock_crossing_bridge_m1_granted_system_tick_s1,
                                    clock_crossing_bridge_m1_qualified_request_system_tick_s1,
                                    clock_crossing_bridge_m1_read_data_valid_system_tick_s1,
                                    clock_crossing_bridge_m1_requests_system_tick_s1,
                                    d1_system_tick_s1_end_xfer,
                                    system_tick_s1_address,
                                    system_tick_s1_chipselect,
                                    system_tick_s1_irq_from_sa,
                                    system_tick_s1_readdata_from_sa,
                                    system_tick_s1_reset_n,
                                    system_tick_s1_write_n,
                                    system_tick_s1_writedata
                                 )
;

  output           clock_crossing_bridge_m1_granted_system_tick_s1;
  output           clock_crossing_bridge_m1_qualified_request_system_tick_s1;
  output           clock_crossing_bridge_m1_read_data_valid_system_tick_s1;
  output           clock_crossing_bridge_m1_requests_system_tick_s1;
  output           d1_system_tick_s1_end_xfer;
  output  [  2: 0] system_tick_s1_address;
  output           system_tick_s1_chipselect;
  output           system_tick_s1_irq_from_sa;
  output  [ 15: 0] system_tick_s1_readdata_from_sa;
  output           system_tick_s1_reset_n;
  output           system_tick_s1_write_n;
  output  [ 15: 0] system_tick_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input            reset_n;
  input            system_tick_s1_irq;
  input   [ 15: 0] system_tick_s1_readdata;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_system_tick_s1;
  wire             clock_crossing_bridge_m1_qualified_request_system_tick_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_system_tick_s1;
  wire             clock_crossing_bridge_m1_requests_system_tick_s1;
  wire             clock_crossing_bridge_m1_saved_grant_system_tick_s1;
  reg              d1_reasons_to_wait;
  reg              d1_system_tick_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_system_tick_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] system_tick_s1_address;
  wire             system_tick_s1_allgrants;
  wire             system_tick_s1_allow_new_arb_cycle;
  wire             system_tick_s1_any_bursting_master_saved_grant;
  wire             system_tick_s1_any_continuerequest;
  wire             system_tick_s1_arb_counter_enable;
  reg              system_tick_s1_arb_share_counter;
  wire             system_tick_s1_arb_share_counter_next_value;
  wire             system_tick_s1_arb_share_set_values;
  wire             system_tick_s1_beginbursttransfer_internal;
  wire             system_tick_s1_begins_xfer;
  wire             system_tick_s1_chipselect;
  wire             system_tick_s1_end_xfer;
  wire             system_tick_s1_firsttransfer;
  wire             system_tick_s1_grant_vector;
  wire             system_tick_s1_in_a_read_cycle;
  wire             system_tick_s1_in_a_write_cycle;
  wire             system_tick_s1_irq_from_sa;
  wire             system_tick_s1_master_qreq_vector;
  wire             system_tick_s1_non_bursting_master_requests;
  wire    [ 15: 0] system_tick_s1_readdata_from_sa;
  reg              system_tick_s1_reg_firsttransfer;
  wire             system_tick_s1_reset_n;
  reg              system_tick_s1_slavearbiterlockenable;
  wire             system_tick_s1_slavearbiterlockenable2;
  wire             system_tick_s1_unreg_firsttransfer;
  wire             system_tick_s1_waits_for_read;
  wire             system_tick_s1_waits_for_write;
  wire             system_tick_s1_write_n;
  wire    [ 15: 0] system_tick_s1_writedata;
  wire             wait_for_system_tick_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~system_tick_s1_end_xfer;
    end


  assign system_tick_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_system_tick_s1));
  //assign system_tick_s1_readdata_from_sa = system_tick_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign system_tick_s1_readdata_from_sa = system_tick_s1_readdata;

  assign clock_crossing_bridge_m1_requests_system_tick_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 5] , 5'b0} == 11'h0) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //system_tick_s1_arb_share_counter set values, which is an e_mux
  assign system_tick_s1_arb_share_set_values = 1;

  //system_tick_s1_non_bursting_master_requests mux, which is an e_mux
  assign system_tick_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_system_tick_s1;

  //system_tick_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign system_tick_s1_any_bursting_master_saved_grant = 0;

  //system_tick_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign system_tick_s1_arb_share_counter_next_value = system_tick_s1_firsttransfer ? (system_tick_s1_arb_share_set_values - 1) : |system_tick_s1_arb_share_counter ? (system_tick_s1_arb_share_counter - 1) : 0;

  //system_tick_s1_allgrants all slave grants, which is an e_mux
  assign system_tick_s1_allgrants = |system_tick_s1_grant_vector;

  //system_tick_s1_end_xfer assignment, which is an e_assign
  assign system_tick_s1_end_xfer = ~(system_tick_s1_waits_for_read | system_tick_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_system_tick_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_system_tick_s1 = system_tick_s1_end_xfer & (~system_tick_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //system_tick_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign system_tick_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_system_tick_s1 & system_tick_s1_allgrants) | (end_xfer_arb_share_counter_term_system_tick_s1 & ~system_tick_s1_non_bursting_master_requests);

  //system_tick_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          system_tick_s1_arb_share_counter <= 0;
      else if (system_tick_s1_arb_counter_enable)
          system_tick_s1_arb_share_counter <= system_tick_s1_arb_share_counter_next_value;
    end


  //system_tick_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          system_tick_s1_slavearbiterlockenable <= 0;
      else if ((|system_tick_s1_master_qreq_vector & end_xfer_arb_share_counter_term_system_tick_s1) | (end_xfer_arb_share_counter_term_system_tick_s1 & ~system_tick_s1_non_bursting_master_requests))
          system_tick_s1_slavearbiterlockenable <= |system_tick_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 system_tick/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = system_tick_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //system_tick_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign system_tick_s1_slavearbiterlockenable2 = |system_tick_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 system_tick/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = system_tick_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //system_tick_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign system_tick_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_system_tick_s1 = clock_crossing_bridge_m1_requests_system_tick_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_system_tick_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_system_tick_s1 = clock_crossing_bridge_m1_granted_system_tick_s1 & clock_crossing_bridge_m1_read & ~system_tick_s1_waits_for_read;

  //system_tick_s1_writedata mux, which is an e_mux
  assign system_tick_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_system_tick_s1 = clock_crossing_bridge_m1_qualified_request_system_tick_s1;

  //clock_crossing_bridge/m1 saved-grant system_tick/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_system_tick_s1 = clock_crossing_bridge_m1_requests_system_tick_s1;

  //allow new arb cycle for system_tick/s1, which is an e_assign
  assign system_tick_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign system_tick_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign system_tick_s1_master_qreq_vector = 1;

  //system_tick_s1_reset_n assignment, which is an e_assign
  assign system_tick_s1_reset_n = reset_n;

  assign system_tick_s1_chipselect = clock_crossing_bridge_m1_granted_system_tick_s1;
  //system_tick_s1_firsttransfer first transaction, which is an e_assign
  assign system_tick_s1_firsttransfer = system_tick_s1_begins_xfer ? system_tick_s1_unreg_firsttransfer : system_tick_s1_reg_firsttransfer;

  //system_tick_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign system_tick_s1_unreg_firsttransfer = ~(system_tick_s1_slavearbiterlockenable & system_tick_s1_any_continuerequest);

  //system_tick_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          system_tick_s1_reg_firsttransfer <= 1'b1;
      else if (system_tick_s1_begins_xfer)
          system_tick_s1_reg_firsttransfer <= system_tick_s1_unreg_firsttransfer;
    end


  //system_tick_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign system_tick_s1_beginbursttransfer_internal = system_tick_s1_begins_xfer;

  //~system_tick_s1_write_n assignment, which is an e_mux
  assign system_tick_s1_write_n = ~(clock_crossing_bridge_m1_granted_system_tick_s1 & clock_crossing_bridge_m1_write);

  //system_tick_s1_address mux, which is an e_mux
  assign system_tick_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_system_tick_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_system_tick_s1_end_xfer <= 1;
      else 
        d1_system_tick_s1_end_xfer <= system_tick_s1_end_xfer;
    end


  //system_tick_s1_waits_for_read in a cycle, which is an e_mux
  assign system_tick_s1_waits_for_read = system_tick_s1_in_a_read_cycle & system_tick_s1_begins_xfer;

  //system_tick_s1_in_a_read_cycle assignment, which is an e_assign
  assign system_tick_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_system_tick_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = system_tick_s1_in_a_read_cycle;

  //system_tick_s1_waits_for_write in a cycle, which is an e_mux
  assign system_tick_s1_waits_for_write = system_tick_s1_in_a_write_cycle & 0;

  //system_tick_s1_in_a_write_cycle assignment, which is an e_assign
  assign system_tick_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_system_tick_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = system_tick_s1_in_a_write_cycle;

  assign wait_for_system_tick_s1_counter = 0;
  //assign system_tick_s1_irq_from_sa = system_tick_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign system_tick_s1_irq_from_sa = system_tick_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //system_tick/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module touchPanel_irq_n_s1_arbitrator (
                                        // inputs:
                                         clk,
                                         clock_crossing_bridge_m1_address_to_slave,
                                         clock_crossing_bridge_m1_latency_counter,
                                         clock_crossing_bridge_m1_nativeaddress,
                                         clock_crossing_bridge_m1_read,
                                         clock_crossing_bridge_m1_write,
                                         clock_crossing_bridge_m1_writedata,
                                         reset_n,
                                         touchPanel_irq_n_s1_irq,
                                         touchPanel_irq_n_s1_readdata,

                                        // outputs:
                                         clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1,
                                         clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1,
                                         clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1,
                                         clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1,
                                         d1_touchPanel_irq_n_s1_end_xfer,
                                         touchPanel_irq_n_s1_address,
                                         touchPanel_irq_n_s1_chipselect,
                                         touchPanel_irq_n_s1_irq_from_sa,
                                         touchPanel_irq_n_s1_readdata_from_sa,
                                         touchPanel_irq_n_s1_reset_n,
                                         touchPanel_irq_n_s1_write_n,
                                         touchPanel_irq_n_s1_writedata
                                      )
;

  output           clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1;
  output           clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1;
  output           clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1;
  output           clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1;
  output           d1_touchPanel_irq_n_s1_end_xfer;
  output  [  1: 0] touchPanel_irq_n_s1_address;
  output           touchPanel_irq_n_s1_chipselect;
  output           touchPanel_irq_n_s1_irq_from_sa;
  output  [ 31: 0] touchPanel_irq_n_s1_readdata_from_sa;
  output           touchPanel_irq_n_s1_reset_n;
  output           touchPanel_irq_n_s1_write_n;
  output  [ 31: 0] touchPanel_irq_n_s1_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input            reset_n;
  input            touchPanel_irq_n_s1_irq;
  input   [ 31: 0] touchPanel_irq_n_s1_readdata;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_saved_grant_touchPanel_irq_n_s1;
  reg              d1_reasons_to_wait;
  reg              d1_touchPanel_irq_n_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_touchPanel_irq_n_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] touchPanel_irq_n_s1_address;
  wire             touchPanel_irq_n_s1_allgrants;
  wire             touchPanel_irq_n_s1_allow_new_arb_cycle;
  wire             touchPanel_irq_n_s1_any_bursting_master_saved_grant;
  wire             touchPanel_irq_n_s1_any_continuerequest;
  wire             touchPanel_irq_n_s1_arb_counter_enable;
  reg              touchPanel_irq_n_s1_arb_share_counter;
  wire             touchPanel_irq_n_s1_arb_share_counter_next_value;
  wire             touchPanel_irq_n_s1_arb_share_set_values;
  wire             touchPanel_irq_n_s1_beginbursttransfer_internal;
  wire             touchPanel_irq_n_s1_begins_xfer;
  wire             touchPanel_irq_n_s1_chipselect;
  wire             touchPanel_irq_n_s1_end_xfer;
  wire             touchPanel_irq_n_s1_firsttransfer;
  wire             touchPanel_irq_n_s1_grant_vector;
  wire             touchPanel_irq_n_s1_in_a_read_cycle;
  wire             touchPanel_irq_n_s1_in_a_write_cycle;
  wire             touchPanel_irq_n_s1_irq_from_sa;
  wire             touchPanel_irq_n_s1_master_qreq_vector;
  wire             touchPanel_irq_n_s1_non_bursting_master_requests;
  wire    [ 31: 0] touchPanel_irq_n_s1_readdata_from_sa;
  reg              touchPanel_irq_n_s1_reg_firsttransfer;
  wire             touchPanel_irq_n_s1_reset_n;
  reg              touchPanel_irq_n_s1_slavearbiterlockenable;
  wire             touchPanel_irq_n_s1_slavearbiterlockenable2;
  wire             touchPanel_irq_n_s1_unreg_firsttransfer;
  wire             touchPanel_irq_n_s1_waits_for_read;
  wire             touchPanel_irq_n_s1_waits_for_write;
  wire             touchPanel_irq_n_s1_write_n;
  wire    [ 31: 0] touchPanel_irq_n_s1_writedata;
  wire             wait_for_touchPanel_irq_n_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~touchPanel_irq_n_s1_end_xfer;
    end


  assign touchPanel_irq_n_s1_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1));
  //assign touchPanel_irq_n_s1_readdata_from_sa = touchPanel_irq_n_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_irq_n_s1_readdata_from_sa = touchPanel_irq_n_s1_readdata;

  assign clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1 = ({clock_crossing_bridge_m1_address_to_slave[10 : 4] , 4'b0} == 11'h280) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //touchPanel_irq_n_s1_arb_share_counter set values, which is an e_mux
  assign touchPanel_irq_n_s1_arb_share_set_values = 1;

  //touchPanel_irq_n_s1_non_bursting_master_requests mux, which is an e_mux
  assign touchPanel_irq_n_s1_non_bursting_master_requests = clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1;

  //touchPanel_irq_n_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign touchPanel_irq_n_s1_any_bursting_master_saved_grant = 0;

  //touchPanel_irq_n_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign touchPanel_irq_n_s1_arb_share_counter_next_value = touchPanel_irq_n_s1_firsttransfer ? (touchPanel_irq_n_s1_arb_share_set_values - 1) : |touchPanel_irq_n_s1_arb_share_counter ? (touchPanel_irq_n_s1_arb_share_counter - 1) : 0;

  //touchPanel_irq_n_s1_allgrants all slave grants, which is an e_mux
  assign touchPanel_irq_n_s1_allgrants = |touchPanel_irq_n_s1_grant_vector;

  //touchPanel_irq_n_s1_end_xfer assignment, which is an e_assign
  assign touchPanel_irq_n_s1_end_xfer = ~(touchPanel_irq_n_s1_waits_for_read | touchPanel_irq_n_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_touchPanel_irq_n_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_touchPanel_irq_n_s1 = touchPanel_irq_n_s1_end_xfer & (~touchPanel_irq_n_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //touchPanel_irq_n_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign touchPanel_irq_n_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_touchPanel_irq_n_s1 & touchPanel_irq_n_s1_allgrants) | (end_xfer_arb_share_counter_term_touchPanel_irq_n_s1 & ~touchPanel_irq_n_s1_non_bursting_master_requests);

  //touchPanel_irq_n_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          touchPanel_irq_n_s1_arb_share_counter <= 0;
      else if (touchPanel_irq_n_s1_arb_counter_enable)
          touchPanel_irq_n_s1_arb_share_counter <= touchPanel_irq_n_s1_arb_share_counter_next_value;
    end


  //touchPanel_irq_n_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          touchPanel_irq_n_s1_slavearbiterlockenable <= 0;
      else if ((|touchPanel_irq_n_s1_master_qreq_vector & end_xfer_arb_share_counter_term_touchPanel_irq_n_s1) | (end_xfer_arb_share_counter_term_touchPanel_irq_n_s1 & ~touchPanel_irq_n_s1_non_bursting_master_requests))
          touchPanel_irq_n_s1_slavearbiterlockenable <= |touchPanel_irq_n_s1_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 touchPanel_irq_n/s1 arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = touchPanel_irq_n_s1_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //touchPanel_irq_n_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign touchPanel_irq_n_s1_slavearbiterlockenable2 = |touchPanel_irq_n_s1_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 touchPanel_irq_n/s1 arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = touchPanel_irq_n_s1_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //touchPanel_irq_n_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign touchPanel_irq_n_s1_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1 = clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1 & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1 = clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1 & clock_crossing_bridge_m1_read & ~touchPanel_irq_n_s1_waits_for_read;

  //touchPanel_irq_n_s1_writedata mux, which is an e_mux
  assign touchPanel_irq_n_s1_writedata = clock_crossing_bridge_m1_writedata;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1 = clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1;

  //clock_crossing_bridge/m1 saved-grant touchPanel_irq_n/s1, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_touchPanel_irq_n_s1 = clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1;

  //allow new arb cycle for touchPanel_irq_n/s1, which is an e_assign
  assign touchPanel_irq_n_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign touchPanel_irq_n_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign touchPanel_irq_n_s1_master_qreq_vector = 1;

  //touchPanel_irq_n_s1_reset_n assignment, which is an e_assign
  assign touchPanel_irq_n_s1_reset_n = reset_n;

  assign touchPanel_irq_n_s1_chipselect = clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1;
  //touchPanel_irq_n_s1_firsttransfer first transaction, which is an e_assign
  assign touchPanel_irq_n_s1_firsttransfer = touchPanel_irq_n_s1_begins_xfer ? touchPanel_irq_n_s1_unreg_firsttransfer : touchPanel_irq_n_s1_reg_firsttransfer;

  //touchPanel_irq_n_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign touchPanel_irq_n_s1_unreg_firsttransfer = ~(touchPanel_irq_n_s1_slavearbiterlockenable & touchPanel_irq_n_s1_any_continuerequest);

  //touchPanel_irq_n_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          touchPanel_irq_n_s1_reg_firsttransfer <= 1'b1;
      else if (touchPanel_irq_n_s1_begins_xfer)
          touchPanel_irq_n_s1_reg_firsttransfer <= touchPanel_irq_n_s1_unreg_firsttransfer;
    end


  //touchPanel_irq_n_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign touchPanel_irq_n_s1_beginbursttransfer_internal = touchPanel_irq_n_s1_begins_xfer;

  //~touchPanel_irq_n_s1_write_n assignment, which is an e_mux
  assign touchPanel_irq_n_s1_write_n = ~(clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1 & clock_crossing_bridge_m1_write);

  //touchPanel_irq_n_s1_address mux, which is an e_mux
  assign touchPanel_irq_n_s1_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_touchPanel_irq_n_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_touchPanel_irq_n_s1_end_xfer <= 1;
      else 
        d1_touchPanel_irq_n_s1_end_xfer <= touchPanel_irq_n_s1_end_xfer;
    end


  //touchPanel_irq_n_s1_waits_for_read in a cycle, which is an e_mux
  assign touchPanel_irq_n_s1_waits_for_read = touchPanel_irq_n_s1_in_a_read_cycle & touchPanel_irq_n_s1_begins_xfer;

  //touchPanel_irq_n_s1_in_a_read_cycle assignment, which is an e_assign
  assign touchPanel_irq_n_s1_in_a_read_cycle = clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1 & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = touchPanel_irq_n_s1_in_a_read_cycle;

  //touchPanel_irq_n_s1_waits_for_write in a cycle, which is an e_mux
  assign touchPanel_irq_n_s1_waits_for_write = touchPanel_irq_n_s1_in_a_write_cycle & 0;

  //touchPanel_irq_n_s1_in_a_write_cycle assignment, which is an e_assign
  assign touchPanel_irq_n_s1_in_a_write_cycle = clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1 & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = touchPanel_irq_n_s1_in_a_write_cycle;

  assign wait_for_touchPanel_irq_n_s1_counter = 0;
  //assign touchPanel_irq_n_s1_irq_from_sa = touchPanel_irq_n_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_irq_n_s1_irq_from_sa = touchPanel_irq_n_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //touchPanel_irq_n/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module touchPanel_spi_spi_control_port_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     clock_crossing_bridge_m1_address_to_slave,
                                                     clock_crossing_bridge_m1_latency_counter,
                                                     clock_crossing_bridge_m1_nativeaddress,
                                                     clock_crossing_bridge_m1_read,
                                                     clock_crossing_bridge_m1_write,
                                                     clock_crossing_bridge_m1_writedata,
                                                     reset_n,
                                                     touchPanel_spi_spi_control_port_dataavailable,
                                                     touchPanel_spi_spi_control_port_endofpacket,
                                                     touchPanel_spi_spi_control_port_irq,
                                                     touchPanel_spi_spi_control_port_readdata,
                                                     touchPanel_spi_spi_control_port_readyfordata,

                                                    // outputs:
                                                     clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port,
                                                     clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port,
                                                     clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port,
                                                     clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port,
                                                     d1_touchPanel_spi_spi_control_port_end_xfer,
                                                     touchPanel_spi_spi_control_port_address,
                                                     touchPanel_spi_spi_control_port_chipselect,
                                                     touchPanel_spi_spi_control_port_dataavailable_from_sa,
                                                     touchPanel_spi_spi_control_port_endofpacket_from_sa,
                                                     touchPanel_spi_spi_control_port_irq_from_sa,
                                                     touchPanel_spi_spi_control_port_read_n,
                                                     touchPanel_spi_spi_control_port_readdata_from_sa,
                                                     touchPanel_spi_spi_control_port_readyfordata_from_sa,
                                                     touchPanel_spi_spi_control_port_reset_n,
                                                     touchPanel_spi_spi_control_port_write_n,
                                                     touchPanel_spi_spi_control_port_writedata
                                                  )
;

  output           clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port;
  output           clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port;
  output           clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port;
  output           clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port;
  output           d1_touchPanel_spi_spi_control_port_end_xfer;
  output  [  2: 0] touchPanel_spi_spi_control_port_address;
  output           touchPanel_spi_spi_control_port_chipselect;
  output           touchPanel_spi_spi_control_port_dataavailable_from_sa;
  output           touchPanel_spi_spi_control_port_endofpacket_from_sa;
  output           touchPanel_spi_spi_control_port_irq_from_sa;
  output           touchPanel_spi_spi_control_port_read_n;
  output  [ 15: 0] touchPanel_spi_spi_control_port_readdata_from_sa;
  output           touchPanel_spi_spi_control_port_readyfordata_from_sa;
  output           touchPanel_spi_spi_control_port_reset_n;
  output           touchPanel_spi_spi_control_port_write_n;
  output  [ 15: 0] touchPanel_spi_spi_control_port_writedata;
  input            clk;
  input   [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  input            clock_crossing_bridge_m1_latency_counter;
  input   [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  input            clock_crossing_bridge_m1_read;
  input            clock_crossing_bridge_m1_write;
  input   [ 31: 0] clock_crossing_bridge_m1_writedata;
  input            reset_n;
  input            touchPanel_spi_spi_control_port_dataavailable;
  input            touchPanel_spi_spi_control_port_endofpacket;
  input            touchPanel_spi_spi_control_port_irq;
  input   [ 15: 0] touchPanel_spi_spi_control_port_readdata;
  input            touchPanel_spi_spi_control_port_readyfordata;

  wire             clock_crossing_bridge_m1_arbiterlock;
  wire             clock_crossing_bridge_m1_arbiterlock2;
  wire             clock_crossing_bridge_m1_continuerequest;
  wire             clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_saved_grant_touchPanel_spi_spi_control_port;
  reg              d1_reasons_to_wait;
  reg              d1_touchPanel_spi_spi_control_port_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] touchPanel_spi_spi_control_port_address;
  wire             touchPanel_spi_spi_control_port_allgrants;
  wire             touchPanel_spi_spi_control_port_allow_new_arb_cycle;
  wire             touchPanel_spi_spi_control_port_any_bursting_master_saved_grant;
  wire             touchPanel_spi_spi_control_port_any_continuerequest;
  wire             touchPanel_spi_spi_control_port_arb_counter_enable;
  reg              touchPanel_spi_spi_control_port_arb_share_counter;
  wire             touchPanel_spi_spi_control_port_arb_share_counter_next_value;
  wire             touchPanel_spi_spi_control_port_arb_share_set_values;
  wire             touchPanel_spi_spi_control_port_beginbursttransfer_internal;
  wire             touchPanel_spi_spi_control_port_begins_xfer;
  wire             touchPanel_spi_spi_control_port_chipselect;
  wire             touchPanel_spi_spi_control_port_dataavailable_from_sa;
  wire             touchPanel_spi_spi_control_port_end_xfer;
  wire             touchPanel_spi_spi_control_port_endofpacket_from_sa;
  wire             touchPanel_spi_spi_control_port_firsttransfer;
  wire             touchPanel_spi_spi_control_port_grant_vector;
  wire             touchPanel_spi_spi_control_port_in_a_read_cycle;
  wire             touchPanel_spi_spi_control_port_in_a_write_cycle;
  wire             touchPanel_spi_spi_control_port_irq_from_sa;
  wire             touchPanel_spi_spi_control_port_master_qreq_vector;
  wire             touchPanel_spi_spi_control_port_non_bursting_master_requests;
  wire             touchPanel_spi_spi_control_port_read_n;
  wire    [ 15: 0] touchPanel_spi_spi_control_port_readdata_from_sa;
  wire             touchPanel_spi_spi_control_port_readyfordata_from_sa;
  reg              touchPanel_spi_spi_control_port_reg_firsttransfer;
  wire             touchPanel_spi_spi_control_port_reset_n;
  reg              touchPanel_spi_spi_control_port_slavearbiterlockenable;
  wire             touchPanel_spi_spi_control_port_slavearbiterlockenable2;
  wire             touchPanel_spi_spi_control_port_unreg_firsttransfer;
  wire             touchPanel_spi_spi_control_port_waits_for_read;
  wire             touchPanel_spi_spi_control_port_waits_for_write;
  wire             touchPanel_spi_spi_control_port_write_n;
  wire    [ 15: 0] touchPanel_spi_spi_control_port_writedata;
  wire             wait_for_touchPanel_spi_spi_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~touchPanel_spi_spi_control_port_end_xfer;
    end


  assign touchPanel_spi_spi_control_port_begins_xfer = ~d1_reasons_to_wait & ((clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port));
  //assign touchPanel_spi_spi_control_port_readdata_from_sa = touchPanel_spi_spi_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_spi_spi_control_port_readdata_from_sa = touchPanel_spi_spi_control_port_readdata;

  assign clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port = ({clock_crossing_bridge_m1_address_to_slave[10 : 5] , 5'b0} == 11'h100) & (clock_crossing_bridge_m1_read | clock_crossing_bridge_m1_write);
  //assign touchPanel_spi_spi_control_port_dataavailable_from_sa = touchPanel_spi_spi_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_spi_spi_control_port_dataavailable_from_sa = touchPanel_spi_spi_control_port_dataavailable;

  //assign touchPanel_spi_spi_control_port_readyfordata_from_sa = touchPanel_spi_spi_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_spi_spi_control_port_readyfordata_from_sa = touchPanel_spi_spi_control_port_readyfordata;

  //touchPanel_spi_spi_control_port_arb_share_counter set values, which is an e_mux
  assign touchPanel_spi_spi_control_port_arb_share_set_values = 1;

  //touchPanel_spi_spi_control_port_non_bursting_master_requests mux, which is an e_mux
  assign touchPanel_spi_spi_control_port_non_bursting_master_requests = clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port;

  //touchPanel_spi_spi_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign touchPanel_spi_spi_control_port_any_bursting_master_saved_grant = 0;

  //touchPanel_spi_spi_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign touchPanel_spi_spi_control_port_arb_share_counter_next_value = touchPanel_spi_spi_control_port_firsttransfer ? (touchPanel_spi_spi_control_port_arb_share_set_values - 1) : |touchPanel_spi_spi_control_port_arb_share_counter ? (touchPanel_spi_spi_control_port_arb_share_counter - 1) : 0;

  //touchPanel_spi_spi_control_port_allgrants all slave grants, which is an e_mux
  assign touchPanel_spi_spi_control_port_allgrants = |touchPanel_spi_spi_control_port_grant_vector;

  //touchPanel_spi_spi_control_port_end_xfer assignment, which is an e_assign
  assign touchPanel_spi_spi_control_port_end_xfer = ~(touchPanel_spi_spi_control_port_waits_for_read | touchPanel_spi_spi_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port = touchPanel_spi_spi_control_port_end_xfer & (~touchPanel_spi_spi_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //touchPanel_spi_spi_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign touchPanel_spi_spi_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port & touchPanel_spi_spi_control_port_allgrants) | (end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port & ~touchPanel_spi_spi_control_port_non_bursting_master_requests);

  //touchPanel_spi_spi_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          touchPanel_spi_spi_control_port_arb_share_counter <= 0;
      else if (touchPanel_spi_spi_control_port_arb_counter_enable)
          touchPanel_spi_spi_control_port_arb_share_counter <= touchPanel_spi_spi_control_port_arb_share_counter_next_value;
    end


  //touchPanel_spi_spi_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          touchPanel_spi_spi_control_port_slavearbiterlockenable <= 0;
      else if ((|touchPanel_spi_spi_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port) | (end_xfer_arb_share_counter_term_touchPanel_spi_spi_control_port & ~touchPanel_spi_spi_control_port_non_bursting_master_requests))
          touchPanel_spi_spi_control_port_slavearbiterlockenable <= |touchPanel_spi_spi_control_port_arb_share_counter_next_value;
    end


  //clock_crossing_bridge/m1 touchPanel_spi/spi_control_port arbiterlock, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock = touchPanel_spi_spi_control_port_slavearbiterlockenable & clock_crossing_bridge_m1_continuerequest;

  //touchPanel_spi_spi_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign touchPanel_spi_spi_control_port_slavearbiterlockenable2 = |touchPanel_spi_spi_control_port_arb_share_counter_next_value;

  //clock_crossing_bridge/m1 touchPanel_spi/spi_control_port arbiterlock2, which is an e_assign
  assign clock_crossing_bridge_m1_arbiterlock2 = touchPanel_spi_spi_control_port_slavearbiterlockenable2 & clock_crossing_bridge_m1_continuerequest;

  //touchPanel_spi_spi_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  assign touchPanel_spi_spi_control_port_any_continuerequest = 1;

  //clock_crossing_bridge_m1_continuerequest continued request, which is an e_assign
  assign clock_crossing_bridge_m1_continuerequest = 1;

  assign clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port = clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port & ~((clock_crossing_bridge_m1_read & ((clock_crossing_bridge_m1_latency_counter != 0))));
  //local readdatavalid clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port, which is an e_mux
  assign clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port = clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port & clock_crossing_bridge_m1_read & ~touchPanel_spi_spi_control_port_waits_for_read;

  //touchPanel_spi_spi_control_port_writedata mux, which is an e_mux
  assign touchPanel_spi_spi_control_port_writedata = clock_crossing_bridge_m1_writedata;

  //assign touchPanel_spi_spi_control_port_endofpacket_from_sa = touchPanel_spi_spi_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_spi_spi_control_port_endofpacket_from_sa = touchPanel_spi_spi_control_port_endofpacket;

  //master is always granted when requested
  assign clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port = clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port;

  //clock_crossing_bridge/m1 saved-grant touchPanel_spi/spi_control_port, which is an e_assign
  assign clock_crossing_bridge_m1_saved_grant_touchPanel_spi_spi_control_port = clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port;

  //allow new arb cycle for touchPanel_spi/spi_control_port, which is an e_assign
  assign touchPanel_spi_spi_control_port_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign touchPanel_spi_spi_control_port_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign touchPanel_spi_spi_control_port_master_qreq_vector = 1;

  //touchPanel_spi_spi_control_port_reset_n assignment, which is an e_assign
  assign touchPanel_spi_spi_control_port_reset_n = reset_n;

  assign touchPanel_spi_spi_control_port_chipselect = clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port;
  //touchPanel_spi_spi_control_port_firsttransfer first transaction, which is an e_assign
  assign touchPanel_spi_spi_control_port_firsttransfer = touchPanel_spi_spi_control_port_begins_xfer ? touchPanel_spi_spi_control_port_unreg_firsttransfer : touchPanel_spi_spi_control_port_reg_firsttransfer;

  //touchPanel_spi_spi_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign touchPanel_spi_spi_control_port_unreg_firsttransfer = ~(touchPanel_spi_spi_control_port_slavearbiterlockenable & touchPanel_spi_spi_control_port_any_continuerequest);

  //touchPanel_spi_spi_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          touchPanel_spi_spi_control_port_reg_firsttransfer <= 1'b1;
      else if (touchPanel_spi_spi_control_port_begins_xfer)
          touchPanel_spi_spi_control_port_reg_firsttransfer <= touchPanel_spi_spi_control_port_unreg_firsttransfer;
    end


  //touchPanel_spi_spi_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign touchPanel_spi_spi_control_port_beginbursttransfer_internal = touchPanel_spi_spi_control_port_begins_xfer;

  //~touchPanel_spi_spi_control_port_read_n assignment, which is an e_mux
  assign touchPanel_spi_spi_control_port_read_n = ~(clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port & clock_crossing_bridge_m1_read);

  //~touchPanel_spi_spi_control_port_write_n assignment, which is an e_mux
  assign touchPanel_spi_spi_control_port_write_n = ~(clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port & clock_crossing_bridge_m1_write);

  //touchPanel_spi_spi_control_port_address mux, which is an e_mux
  assign touchPanel_spi_spi_control_port_address = clock_crossing_bridge_m1_nativeaddress;

  //d1_touchPanel_spi_spi_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_touchPanel_spi_spi_control_port_end_xfer <= 1;
      else 
        d1_touchPanel_spi_spi_control_port_end_xfer <= touchPanel_spi_spi_control_port_end_xfer;
    end


  //touchPanel_spi_spi_control_port_waits_for_read in a cycle, which is an e_mux
  assign touchPanel_spi_spi_control_port_waits_for_read = touchPanel_spi_spi_control_port_in_a_read_cycle & touchPanel_spi_spi_control_port_begins_xfer;

  //touchPanel_spi_spi_control_port_in_a_read_cycle assignment, which is an e_assign
  assign touchPanel_spi_spi_control_port_in_a_read_cycle = clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port & clock_crossing_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = touchPanel_spi_spi_control_port_in_a_read_cycle;

  //touchPanel_spi_spi_control_port_waits_for_write in a cycle, which is an e_mux
  assign touchPanel_spi_spi_control_port_waits_for_write = touchPanel_spi_spi_control_port_in_a_write_cycle & touchPanel_spi_spi_control_port_begins_xfer;

  //touchPanel_spi_spi_control_port_in_a_write_cycle assignment, which is an e_assign
  assign touchPanel_spi_spi_control_port_in_a_write_cycle = clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port & clock_crossing_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = touchPanel_spi_spi_control_port_in_a_write_cycle;

  assign wait_for_touchPanel_spi_spi_control_port_counter = 0;
  //assign touchPanel_spi_spi_control_port_irq_from_sa = touchPanel_spi_spi_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign touchPanel_spi_spi_control_port_irq_from_sa = touchPanel_spi_spi_control_port_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //touchPanel_spi/spi_control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tristate_bridge_avalon_slave_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  flash_ssram_pipeline_bridge_m1_address_to_slave,
                                                  flash_ssram_pipeline_bridge_m1_burstcount,
                                                  flash_ssram_pipeline_bridge_m1_byteenable,
                                                  flash_ssram_pipeline_bridge_m1_chipselect,
                                                  flash_ssram_pipeline_bridge_m1_dbs_address,
                                                  flash_ssram_pipeline_bridge_m1_dbs_write_16,
                                                  flash_ssram_pipeline_bridge_m1_dbs_write_32,
                                                  flash_ssram_pipeline_bridge_m1_latency_counter,
                                                  flash_ssram_pipeline_bridge_m1_read,
                                                  flash_ssram_pipeline_bridge_m1_write,
                                                  reset_n,

                                                 // outputs:
                                                  adsc_n_to_the_ssram,
                                                  bw_n_to_the_ssram,
                                                  bwe_n_to_the_ssram,
                                                  chipenable1_n_to_the_ssram,
                                                  d1_tristate_bridge_avalon_slave_end_xfer,
                                                  flash_s1_wait_counter_eq_0,
                                                  flash_ssram_pipeline_bridge_m1_byteenable_flash_s1,
                                                  flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1,
                                                  flash_ssram_pipeline_bridge_m1_granted_flash_s1,
                                                  flash_ssram_pipeline_bridge_m1_granted_ssram_s1,
                                                  flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1,
                                                  flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1,
                                                  flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1,
                                                  flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1,
                                                  flash_ssram_pipeline_bridge_m1_requests_flash_s1,
                                                  flash_ssram_pipeline_bridge_m1_requests_ssram_s1,
                                                  incoming_tristate_bridge_data,
                                                  incoming_tristate_bridge_data_with_Xs_converted_to_0,
                                                  outputenable_n_to_the_ssram,
                                                  read_n_to_the_flash,
                                                  reset_n_to_the_ssram,
                                                  select_n_to_the_flash,
                                                  tristate_bridge_address,
                                                  tristate_bridge_data,
                                                  write_n_to_the_flash
                                               )
;

  output           adsc_n_to_the_ssram;
  output  [  3: 0] bw_n_to_the_ssram;
  output           bwe_n_to_the_ssram;
  output           chipenable1_n_to_the_ssram;
  output           d1_tristate_bridge_avalon_slave_end_xfer;
  output           flash_s1_wait_counter_eq_0;
  output  [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1;
  output  [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1;
  output           flash_ssram_pipeline_bridge_m1_granted_flash_s1;
  output           flash_ssram_pipeline_bridge_m1_granted_ssram_s1;
  output           flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1;
  output           flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1;
  output           flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1;
  output           flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1;
  output           flash_ssram_pipeline_bridge_m1_requests_flash_s1;
  output           flash_ssram_pipeline_bridge_m1_requests_ssram_s1;
  output  [ 31: 0] incoming_tristate_bridge_data;
  output  [ 15: 0] incoming_tristate_bridge_data_with_Xs_converted_to_0;
  output           outputenable_n_to_the_ssram;
  output           read_n_to_the_flash;
  output           reset_n_to_the_ssram;
  output           select_n_to_the_flash;
  output  [ 23: 0] tristate_bridge_address;
  inout   [ 31: 0] tristate_bridge_data;
  output           write_n_to_the_flash;
  input            clk;
  input   [ 24: 0] flash_ssram_pipeline_bridge_m1_address_to_slave;
  input            flash_ssram_pipeline_bridge_m1_burstcount;
  input   [ 31: 0] flash_ssram_pipeline_bridge_m1_byteenable;
  input            flash_ssram_pipeline_bridge_m1_chipselect;
  input   [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_address;
  input   [ 15: 0] flash_ssram_pipeline_bridge_m1_dbs_write_16;
  input   [ 31: 0] flash_ssram_pipeline_bridge_m1_dbs_write_32;
  input   [  2: 0] flash_ssram_pipeline_bridge_m1_latency_counter;
  input            flash_ssram_pipeline_bridge_m1_read;
  input            flash_ssram_pipeline_bridge_m1_write;
  input            reset_n;

  reg              adsc_n_to_the_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg     [  3: 0] bw_n_to_the_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              bwe_n_to_the_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              chipenable1_n_to_the_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [ 31: 0] d1_outgoing_tristate_bridge_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              d1_tristate_bridge_avalon_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave;
  wire    [  3: 0] flash_s1_counter_load_value;
  wire             flash_s1_in_a_read_cycle;
  wire             flash_s1_in_a_write_cycle;
  reg     [  3: 0] flash_s1_wait_counter;
  wire             flash_s1_wait_counter_eq_0;
  wire             flash_s1_waits_for_read;
  wire             flash_s1_waits_for_write;
  wire             flash_s1_with_write_latency;
  wire             flash_ssram_pipeline_bridge_m1_arbiterlock;
  wire             flash_ssram_pipeline_bridge_m1_arbiterlock2;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_0;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_1;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_10;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_11;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_12;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_13;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_14;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_15;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_2;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_3;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_4;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_5;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_6;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_7;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_8;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_9;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_0;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_1;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_2;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_3;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_4;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_5;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_6;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_7;
  wire             flash_ssram_pipeline_bridge_m1_continuerequest;
  wire             flash_ssram_pipeline_bridge_m1_granted_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_granted_ssram_s1;
  wire             flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1;
  wire             flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1;
  reg     [  1: 0] flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register;
  wire             flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register_in;
  wire             flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1;
  reg     [  3: 0] flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register;
  wire             flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register_in;
  wire             flash_ssram_pipeline_bridge_m1_requests_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_requests_ssram_s1;
  wire             flash_ssram_pipeline_bridge_m1_saved_grant_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_saved_grant_ssram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 31: 0] incoming_tristate_bridge_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  wire             incoming_tristate_bridge_data_bit_0_is_x;
  wire             incoming_tristate_bridge_data_bit_10_is_x;
  wire             incoming_tristate_bridge_data_bit_11_is_x;
  wire             incoming_tristate_bridge_data_bit_12_is_x;
  wire             incoming_tristate_bridge_data_bit_13_is_x;
  wire             incoming_tristate_bridge_data_bit_14_is_x;
  wire             incoming_tristate_bridge_data_bit_15_is_x;
  wire             incoming_tristate_bridge_data_bit_1_is_x;
  wire             incoming_tristate_bridge_data_bit_2_is_x;
  wire             incoming_tristate_bridge_data_bit_3_is_x;
  wire             incoming_tristate_bridge_data_bit_4_is_x;
  wire             incoming_tristate_bridge_data_bit_5_is_x;
  wire             incoming_tristate_bridge_data_bit_6_is_x;
  wire             incoming_tristate_bridge_data_bit_7_is_x;
  wire             incoming_tristate_bridge_data_bit_8_is_x;
  wire             incoming_tristate_bridge_data_bit_9_is_x;
  wire    [ 15: 0] incoming_tristate_bridge_data_with_Xs_converted_to_0;
  wire    [ 31: 0] outgoing_tristate_bridge_data;
  reg              outputenable_n_to_the_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             p1_adsc_n_to_the_ssram;
  wire    [  3: 0] p1_bw_n_to_the_ssram;
  wire             p1_bwe_n_to_the_ssram;
  wire             p1_chipenable1_n_to_the_ssram;
  wire    [  1: 0] p1_flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register;
  wire    [  3: 0] p1_flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register;
  wire             p1_outputenable_n_to_the_ssram;
  wire             p1_read_n_to_the_flash;
  wire             p1_reset_n_to_the_ssram;
  wire             p1_select_n_to_the_flash;
  wire    [ 23: 0] p1_tristate_bridge_address;
  wire             p1_write_n_to_the_flash;
  reg              read_n_to_the_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              reset_n_to_the_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              select_n_to_the_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             ssram_s1_in_a_read_cycle;
  wire             ssram_s1_in_a_write_cycle;
  wire             ssram_s1_waits_for_read;
  wire             ssram_s1_waits_for_write;
  wire             ssram_s1_with_write_latency;
  wire             time_to_write;
  reg     [ 23: 0] tristate_bridge_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             tristate_bridge_avalon_slave_allgrants;
  wire             tristate_bridge_avalon_slave_allow_new_arb_cycle;
  wire             tristate_bridge_avalon_slave_any_bursting_master_saved_grant;
  wire             tristate_bridge_avalon_slave_any_continuerequest;
  wire             tristate_bridge_avalon_slave_arb_counter_enable;
  reg     [  4: 0] tristate_bridge_avalon_slave_arb_share_counter;
  wire    [  4: 0] tristate_bridge_avalon_slave_arb_share_counter_next_value;
  wire    [  4: 0] tristate_bridge_avalon_slave_arb_share_set_values;
  wire             tristate_bridge_avalon_slave_beginbursttransfer_internal;
  wire             tristate_bridge_avalon_slave_begins_xfer;
  wire             tristate_bridge_avalon_slave_end_xfer;
  wire             tristate_bridge_avalon_slave_firsttransfer;
  wire             tristate_bridge_avalon_slave_grant_vector;
  wire             tristate_bridge_avalon_slave_master_qreq_vector;
  wire             tristate_bridge_avalon_slave_non_bursting_master_requests;
  wire             tristate_bridge_avalon_slave_read_pending;
  reg              tristate_bridge_avalon_slave_reg_firsttransfer;
  reg              tristate_bridge_avalon_slave_slavearbiterlockenable;
  wire             tristate_bridge_avalon_slave_slavearbiterlockenable2;
  wire             tristate_bridge_avalon_slave_unreg_firsttransfer;
  wire             tristate_bridge_avalon_slave_write_pending;
  wire    [ 31: 0] tristate_bridge_data;
  wire             wait_for_flash_s1_counter;
  wire             wait_for_ssram_s1_counter;
  reg              write_n_to_the_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tristate_bridge_avalon_slave_end_xfer;
    end


  assign tristate_bridge_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 | flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1));
  assign flash_ssram_pipeline_bridge_m1_requests_flash_s1 = ({flash_ssram_pipeline_bridge_m1_address_to_slave[24] , 24'b0} == 25'h2000000) & flash_ssram_pipeline_bridge_m1_chipselect;
  //~select_n_to_the_flash of type chipselect to ~p1_select_n_to_the_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_flash <= ~0;
      else 
        select_n_to_the_flash <= p1_select_n_to_the_flash;
    end


  //~chipenable1_n_to_the_ssram of type chipselect to ~p1_chipenable1_n_to_the_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          chipenable1_n_to_the_ssram <= ~0;
      else 
        chipenable1_n_to_the_ssram <= p1_chipenable1_n_to_the_ssram;
    end


  assign tristate_bridge_avalon_slave_write_pending = 0;
  //tristate_bridge/avalon_slave read pending calc, which is an e_assign
  assign tristate_bridge_avalon_slave_read_pending = |flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register[1 : 0];

  //tristate_bridge_avalon_slave_arb_share_counter set values, which is an e_mux
  assign tristate_bridge_avalon_slave_arb_share_set_values = (flash_ssram_pipeline_bridge_m1_granted_flash_s1)? 16 :
    (flash_ssram_pipeline_bridge_m1_granted_ssram_s1)? 8 :
    1;

  //tristate_bridge_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign tristate_bridge_avalon_slave_non_bursting_master_requests = flash_ssram_pipeline_bridge_m1_requests_flash_s1 |
    flash_ssram_pipeline_bridge_m1_requests_ssram_s1;

  //tristate_bridge_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign tristate_bridge_avalon_slave_any_bursting_master_saved_grant = 0;

  //tristate_bridge_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign tristate_bridge_avalon_slave_arb_share_counter_next_value = tristate_bridge_avalon_slave_firsttransfer ? (tristate_bridge_avalon_slave_arb_share_set_values - 1) : |tristate_bridge_avalon_slave_arb_share_counter ? (tristate_bridge_avalon_slave_arb_share_counter - 1) : 0;

  //tristate_bridge_avalon_slave_allgrants all slave grants, which is an e_mux
  assign tristate_bridge_avalon_slave_allgrants = (|tristate_bridge_avalon_slave_grant_vector) |
    (|tristate_bridge_avalon_slave_grant_vector);

  //tristate_bridge_avalon_slave_end_xfer assignment, which is an e_assign
  assign tristate_bridge_avalon_slave_end_xfer = ~(flash_s1_waits_for_read | flash_s1_waits_for_write | ssram_s1_waits_for_read | ssram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave = tristate_bridge_avalon_slave_end_xfer & (~tristate_bridge_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tristate_bridge_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign tristate_bridge_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave & tristate_bridge_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave & ~tristate_bridge_avalon_slave_non_bursting_master_requests);

  //tristate_bridge_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tristate_bridge_avalon_slave_arb_share_counter <= 0;
      else if (tristate_bridge_avalon_slave_arb_counter_enable)
          tristate_bridge_avalon_slave_arb_share_counter <= tristate_bridge_avalon_slave_arb_share_counter_next_value;
    end


  //tristate_bridge_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tristate_bridge_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|tristate_bridge_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave) | (end_xfer_arb_share_counter_term_tristate_bridge_avalon_slave & ~tristate_bridge_avalon_slave_non_bursting_master_requests))
          tristate_bridge_avalon_slave_slavearbiterlockenable <= |tristate_bridge_avalon_slave_arb_share_counter_next_value;
    end


  //flash_ssram_pipeline_bridge/m1 tristate_bridge/avalon_slave arbiterlock, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_arbiterlock = tristate_bridge_avalon_slave_slavearbiterlockenable & flash_ssram_pipeline_bridge_m1_continuerequest;

  //tristate_bridge_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tristate_bridge_avalon_slave_slavearbiterlockenable2 = |tristate_bridge_avalon_slave_arb_share_counter_next_value;

  //flash_ssram_pipeline_bridge/m1 tristate_bridge/avalon_slave arbiterlock2, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_arbiterlock2 = tristate_bridge_avalon_slave_slavearbiterlockenable2 & flash_ssram_pipeline_bridge_m1_continuerequest;

  //tristate_bridge_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tristate_bridge_avalon_slave_any_continuerequest = 1;

  //flash_ssram_pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_continuerequest = 1;

  assign flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 = flash_ssram_pipeline_bridge_m1_requests_flash_s1 & ~(((flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & (tristate_bridge_avalon_slave_write_pending | (tristate_bridge_avalon_slave_read_pending) | (2 < flash_ssram_pipeline_bridge_m1_latency_counter))) | ((tristate_bridge_avalon_slave_read_pending | !flash_ssram_pipeline_bridge_m1_byteenable_flash_s1) & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect)));
  //flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register_in = flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & ~flash_s1_waits_for_read;

  //shift register p1 flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register = {flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register, flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register_in};

  //flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register <= p1_flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register;
    end


  //local readdatavalid flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1 = flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1_shift_register[1];

  //tristate_bridge_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_tristate_bridge_data <= 0;
      else 
        incoming_tristate_bridge_data <= tristate_bridge_data;
    end


  //flash_s1_with_write_latency assignment, which is an e_assign
  assign flash_s1_with_write_latency = in_a_write_cycle & (flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (flash_s1_with_write_latency)? 1 :
    (ssram_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_tristate_bridge_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_tristate_bridge_data <= 0;
      else 
        d1_outgoing_tristate_bridge_data <= outgoing_tristate_bridge_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else 
        d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_tristate_bridge_data tristate driver, which is an e_assign
  assign tristate_bridge_data = (d1_in_a_write_cycle)? d1_outgoing_tristate_bridge_data:{32{1'bz}};

  //outgoing_tristate_bridge_data mux, which is an e_mux
  assign outgoing_tristate_bridge_data = (flash_ssram_pipeline_bridge_m1_granted_flash_s1)? flash_ssram_pipeline_bridge_m1_dbs_write_16 :
    flash_ssram_pipeline_bridge_m1_dbs_write_32;

  assign flash_ssram_pipeline_bridge_m1_requests_ssram_s1 = ({flash_ssram_pipeline_bridge_m1_address_to_slave[24 : 20] , 20'b0} == 25'h3000000) & flash_ssram_pipeline_bridge_m1_chipselect;
  assign flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1 = flash_ssram_pipeline_bridge_m1_requests_ssram_s1 & ~(((flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & (tristate_bridge_avalon_slave_write_pending | (tristate_bridge_avalon_slave_read_pending & !((((|flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register[1 : 0]))))) | (4 < flash_ssram_pipeline_bridge_m1_latency_counter))) | ((tristate_bridge_avalon_slave_read_pending | !flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1) & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect)));
  //flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register_in = flash_ssram_pipeline_bridge_m1_granted_ssram_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect) & ~ssram_s1_waits_for_read;

  //shift register p1 flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register = {flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register, flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register_in};

  //flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register <= 0;
      else 
        flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register <= p1_flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register;
    end


  //local readdatavalid flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1, which is an e_mux
  assign flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1 = flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register[3];

  //ssram_s1_with_write_latency assignment, which is an e_assign
  assign ssram_s1_with_write_latency = in_a_write_cycle & (flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1);

  //master is always granted when requested
  assign flash_ssram_pipeline_bridge_m1_granted_flash_s1 = flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1;

  //flash_ssram_pipeline_bridge/m1 saved-grant flash/s1, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_saved_grant_flash_s1 = flash_ssram_pipeline_bridge_m1_requests_flash_s1;

  //allow new arb cycle for tristate_bridge/avalon_slave, which is an e_assign
  assign tristate_bridge_avalon_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tristate_bridge_avalon_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tristate_bridge_avalon_slave_master_qreq_vector = 1;

  //master is always granted when requested
  assign flash_ssram_pipeline_bridge_m1_granted_ssram_s1 = flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1;

  //flash_ssram_pipeline_bridge/m1 saved-grant ssram/s1, which is an e_assign
  assign flash_ssram_pipeline_bridge_m1_saved_grant_ssram_s1 = flash_ssram_pipeline_bridge_m1_requests_ssram_s1;

  assign p1_select_n_to_the_flash = ~flash_ssram_pipeline_bridge_m1_granted_flash_s1;
  //tristate_bridge_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign tristate_bridge_avalon_slave_firsttransfer = tristate_bridge_avalon_slave_begins_xfer ? tristate_bridge_avalon_slave_unreg_firsttransfer : tristate_bridge_avalon_slave_reg_firsttransfer;

  //tristate_bridge_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign tristate_bridge_avalon_slave_unreg_firsttransfer = ~(tristate_bridge_avalon_slave_slavearbiterlockenable & tristate_bridge_avalon_slave_any_continuerequest);

  //tristate_bridge_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tristate_bridge_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (tristate_bridge_avalon_slave_begins_xfer)
          tristate_bridge_avalon_slave_reg_firsttransfer <= tristate_bridge_avalon_slave_unreg_firsttransfer;
    end


  //tristate_bridge_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tristate_bridge_avalon_slave_beginbursttransfer_internal = tristate_bridge_avalon_slave_begins_xfer;

  //~read_n_to_the_flash of type read to ~p1_read_n_to_the_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_n_to_the_flash <= ~0;
      else 
        read_n_to_the_flash <= p1_read_n_to_the_flash;
    end


  //~p1_read_n_to_the_flash assignment, which is an e_mux
  assign p1_read_n_to_the_flash = ~(((flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect)))& ~tristate_bridge_avalon_slave_begins_xfer & (flash_s1_wait_counter < 7));

  //~write_n_to_the_flash of type write to ~p1_write_n_to_the_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_n_to_the_flash <= ~0;
      else 
        write_n_to_the_flash <= p1_write_n_to_the_flash;
    end


  //~p1_write_n_to_the_flash assignment, which is an e_mux
  assign p1_write_n_to_the_flash = ~(((flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect))) & ~tristate_bridge_avalon_slave_begins_xfer & (flash_s1_wait_counter >= 2) & (flash_s1_wait_counter < 9));

  //tristate_bridge_address of type address to p1_tristate_bridge_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tristate_bridge_address <= 0;
      else 
        tristate_bridge_address <= p1_tristate_bridge_address;
    end


  //p1_tristate_bridge_address mux, which is an e_mux
  assign p1_tristate_bridge_address = (flash_ssram_pipeline_bridge_m1_granted_flash_s1)? ({flash_ssram_pipeline_bridge_m1_address_to_slave >> 5,
    flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1],
    {1 {1'b0}}}) :
    ({flash_ssram_pipeline_bridge_m1_address_to_slave >> 5,
    flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2],
    {2 {1'b0}}});

  //d1_tristate_bridge_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tristate_bridge_avalon_slave_end_xfer <= 1;
      else 
        d1_tristate_bridge_avalon_slave_end_xfer <= tristate_bridge_avalon_slave_end_xfer;
    end


  //flash_s1_waits_for_read in a cycle, which is an e_mux
  assign flash_s1_waits_for_read = flash_s1_in_a_read_cycle & wait_for_flash_s1_counter;

  //flash_s1_in_a_read_cycle assignment, which is an e_assign
  assign flash_s1_in_a_read_cycle = flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = flash_s1_in_a_read_cycle |
    ssram_s1_in_a_read_cycle;

  //flash_s1_waits_for_write in a cycle, which is an e_mux
  assign flash_s1_waits_for_write = flash_s1_in_a_write_cycle & wait_for_flash_s1_counter;

  //flash_s1_in_a_write_cycle assignment, which is an e_assign
  assign flash_s1_in_a_write_cycle = flash_ssram_pipeline_bridge_m1_granted_flash_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = flash_s1_in_a_write_cycle |
    ssram_s1_in_a_write_cycle;

  assign flash_s1_wait_counter_eq_0 = flash_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_s1_wait_counter <= 0;
      else 
        flash_s1_wait_counter <= flash_s1_counter_load_value;
    end


  assign flash_s1_counter_load_value = ((flash_s1_in_a_read_cycle & tristate_bridge_avalon_slave_begins_xfer))? 8 :
    ((flash_s1_in_a_write_cycle & tristate_bridge_avalon_slave_begins_xfer))? 10 :
    (~flash_s1_wait_counter_eq_0)? flash_s1_wait_counter - 1 :
    0;

  assign wait_for_flash_s1_counter = tristate_bridge_avalon_slave_begins_xfer | ~flash_s1_wait_counter_eq_0;
  assign {flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_15,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_14,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_13,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_12,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_11,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_10,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_9,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_8,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_7,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_6,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_5,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_4,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_3,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_2,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_1,
flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_0} = flash_ssram_pipeline_bridge_m1_byteenable;
  assign flash_ssram_pipeline_bridge_m1_byteenable_flash_s1 = ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 0))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_0 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 1))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_1 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 2))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_2 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 3))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_3 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 4))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_4 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 5))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_5 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 6))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_6 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 7))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_7 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 8))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_8 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 9))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_9 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 10))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_10 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 11))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_11 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 12))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_12 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 13))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_13 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 1] == 14))? flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_14 :
    flash_ssram_pipeline_bridge_m1_byteenable_flash_s1_segment_15;

  //~adsc_n_to_the_ssram of type begintransfer to ~p1_adsc_n_to_the_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          adsc_n_to_the_ssram <= ~0;
      else 
        adsc_n_to_the_ssram <= p1_adsc_n_to_the_ssram;
    end


  assign p1_adsc_n_to_the_ssram = ~tristate_bridge_avalon_slave_begins_xfer;
  //~outputenable_n_to_the_ssram of type outputenable to ~p1_outputenable_n_to_the_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          outputenable_n_to_the_ssram <= ~0;
      else 
        outputenable_n_to_the_ssram <= p1_outputenable_n_to_the_ssram;
    end


  //~p1_outputenable_n_to_the_ssram assignment, which is an e_mux
  assign p1_outputenable_n_to_the_ssram = ~((|flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register[1 : 0]) | ssram_s1_in_a_read_cycle);

  //reset_n_to_the_ssram of type reset_n to p1_reset_n_to_the_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reset_n_to_the_ssram <= 0;
      else 
        reset_n_to_the_ssram <= p1_reset_n_to_the_ssram;
    end


  //p1_reset_n_to_the_ssram assignment, which is an e_assign
  assign p1_reset_n_to_the_ssram = reset_n;

  assign p1_chipenable1_n_to_the_ssram = ~(flash_ssram_pipeline_bridge_m1_granted_ssram_s1 | (|flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1_shift_register[1 : 0]));
  //~bwe_n_to_the_ssram of type write to ~p1_bwe_n_to_the_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          bwe_n_to_the_ssram <= ~0;
      else 
        bwe_n_to_the_ssram <= p1_bwe_n_to_the_ssram;
    end


  //~bw_n_to_the_ssram of type byteenable to ~p1_bw_n_to_the_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          bw_n_to_the_ssram <= ~0;
      else 
        bw_n_to_the_ssram <= p1_bw_n_to_the_ssram;
    end


  //~p1_bwe_n_to_the_ssram assignment, which is an e_mux
  assign p1_bwe_n_to_the_ssram = ~(flash_ssram_pipeline_bridge_m1_granted_ssram_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect));

  //ssram_s1_waits_for_read in a cycle, which is an e_mux
  assign ssram_s1_waits_for_read = ssram_s1_in_a_read_cycle & 0;

  //ssram_s1_in_a_read_cycle assignment, which is an e_assign
  assign ssram_s1_in_a_read_cycle = flash_ssram_pipeline_bridge_m1_granted_ssram_s1 & (flash_ssram_pipeline_bridge_m1_read & flash_ssram_pipeline_bridge_m1_chipselect);

  //ssram_s1_waits_for_write in a cycle, which is an e_mux
  assign ssram_s1_waits_for_write = ssram_s1_in_a_write_cycle & 0;

  //ssram_s1_in_a_write_cycle assignment, which is an e_assign
  assign ssram_s1_in_a_write_cycle = flash_ssram_pipeline_bridge_m1_granted_ssram_s1 & (flash_ssram_pipeline_bridge_m1_write & flash_ssram_pipeline_bridge_m1_chipselect);

  assign wait_for_ssram_s1_counter = 0;
  //~p1_bw_n_to_the_ssram byte enable port mux, which is an e_mux
  assign p1_bw_n_to_the_ssram = ~((flash_ssram_pipeline_bridge_m1_granted_ssram_s1)? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1 :
    -1);

  assign {flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_7,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_6,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_5,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_4,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_3,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_2,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_1,
flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_0} = flash_ssram_pipeline_bridge_m1_byteenable;
  assign flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1 = ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 0))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_0 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 1))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_1 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 2))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_2 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 3))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_3 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 4))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_4 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 5))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_5 :
    ((flash_ssram_pipeline_bridge_m1_dbs_address[4 : 2] == 6))? flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_6 :
    flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1_segment_7;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //incoming_tristate_bridge_data_bit_0_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_0_is_x = ^(incoming_tristate_bridge_data[0]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[0] = incoming_tristate_bridge_data_bit_0_is_x ? 1'b0 : incoming_tristate_bridge_data[0];

  //incoming_tristate_bridge_data_bit_1_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_1_is_x = ^(incoming_tristate_bridge_data[1]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[1] = incoming_tristate_bridge_data_bit_1_is_x ? 1'b0 : incoming_tristate_bridge_data[1];

  //incoming_tristate_bridge_data_bit_2_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_2_is_x = ^(incoming_tristate_bridge_data[2]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[2] = incoming_tristate_bridge_data_bit_2_is_x ? 1'b0 : incoming_tristate_bridge_data[2];

  //incoming_tristate_bridge_data_bit_3_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_3_is_x = ^(incoming_tristate_bridge_data[3]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[3] = incoming_tristate_bridge_data_bit_3_is_x ? 1'b0 : incoming_tristate_bridge_data[3];

  //incoming_tristate_bridge_data_bit_4_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_4_is_x = ^(incoming_tristate_bridge_data[4]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[4] = incoming_tristate_bridge_data_bit_4_is_x ? 1'b0 : incoming_tristate_bridge_data[4];

  //incoming_tristate_bridge_data_bit_5_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_5_is_x = ^(incoming_tristate_bridge_data[5]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[5] = incoming_tristate_bridge_data_bit_5_is_x ? 1'b0 : incoming_tristate_bridge_data[5];

  //incoming_tristate_bridge_data_bit_6_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_6_is_x = ^(incoming_tristate_bridge_data[6]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[6] = incoming_tristate_bridge_data_bit_6_is_x ? 1'b0 : incoming_tristate_bridge_data[6];

  //incoming_tristate_bridge_data_bit_7_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_7_is_x = ^(incoming_tristate_bridge_data[7]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[7] = incoming_tristate_bridge_data_bit_7_is_x ? 1'b0 : incoming_tristate_bridge_data[7];

  //incoming_tristate_bridge_data_bit_8_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_8_is_x = ^(incoming_tristate_bridge_data[8]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[8] = incoming_tristate_bridge_data_bit_8_is_x ? 1'b0 : incoming_tristate_bridge_data[8];

  //incoming_tristate_bridge_data_bit_9_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_9_is_x = ^(incoming_tristate_bridge_data[9]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[9] = incoming_tristate_bridge_data_bit_9_is_x ? 1'b0 : incoming_tristate_bridge_data[9];

  //incoming_tristate_bridge_data_bit_10_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_10_is_x = ^(incoming_tristate_bridge_data[10]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[10] = incoming_tristate_bridge_data_bit_10_is_x ? 1'b0 : incoming_tristate_bridge_data[10];

  //incoming_tristate_bridge_data_bit_11_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_11_is_x = ^(incoming_tristate_bridge_data[11]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[11] = incoming_tristate_bridge_data_bit_11_is_x ? 1'b0 : incoming_tristate_bridge_data[11];

  //incoming_tristate_bridge_data_bit_12_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_12_is_x = ^(incoming_tristate_bridge_data[12]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[12] = incoming_tristate_bridge_data_bit_12_is_x ? 1'b0 : incoming_tristate_bridge_data[12];

  //incoming_tristate_bridge_data_bit_13_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_13_is_x = ^(incoming_tristate_bridge_data[13]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[13] = incoming_tristate_bridge_data_bit_13_is_x ? 1'b0 : incoming_tristate_bridge_data[13];

  //incoming_tristate_bridge_data_bit_14_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_14_is_x = ^(incoming_tristate_bridge_data[14]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[14] = incoming_tristate_bridge_data_bit_14_is_x ? 1'b0 : incoming_tristate_bridge_data[14];

  //incoming_tristate_bridge_data_bit_15_is_x x check, which is an e_assign_is_x
  assign incoming_tristate_bridge_data_bit_15_is_x = ^(incoming_tristate_bridge_data[15]) === 1'bx;

  //Crush incoming_tristate_bridge_data_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
  assign incoming_tristate_bridge_data_with_Xs_converted_to_0[15] = incoming_tristate_bridge_data_bit_15_is_x ? 1'b0 : incoming_tristate_bridge_data[15];

  //flash/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //flash_ssram_pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (flash_ssram_pipeline_bridge_m1_requests_flash_s1 && (flash_ssram_pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: flash_ssram_pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave flash/s1", $time);
          $stop;
        end
    end


  //ssram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (flash_ssram_pipeline_bridge_m1_granted_flash_s1 + flash_ssram_pipeline_bridge_m1_granted_ssram_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (flash_ssram_pipeline_bridge_m1_saved_grant_flash_s1 + flash_ssram_pipeline_bridge_m1_saved_grant_ssram_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign incoming_tristate_bridge_data_with_Xs_converted_to_0 = incoming_tristate_bridge_data;
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tristate_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_reset_system_clk_domain_synch_module (
                                                     // inputs:
                                                      clk,
                                                      data_in,
                                                      reset_n,

                                                     // outputs:
                                                      data_out
                                                   )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_reset_frame_buffer_phy_clk_out_domain_synch_module (
                                                                   // inputs:
                                                                    clk,
                                                                    data_in,
                                                                    reset_n,

                                                                   // outputs:
                                                                    data_out
                                                                 )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_reset_slow_clk_domain_synch_module (
                                                   // inputs:
                                                    clk,
                                                    data_in,
                                                    reset_n,

                                                   // outputs:
                                                    data_out
                                                 )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system_reset_video_clk_domain_synch_module (
                                                    // inputs:
                                                     clk,
                                                     data_in,
                                                     reset_n,

                                                    // outputs:
                                                     data_out
                                                  )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module system (
                // 1) global signals:
                 ext_clk_one,
                 frame_buffer_aux_full_rate_clk_out,
                 frame_buffer_aux_half_rate_clk_out,
                 frame_buffer_phy_clk_out,
                 reset_n,
                 slow_clk,
                 system_clk,
                 video_clk,

                // the_frame_buffer
                 global_reset_n_to_the_frame_buffer,
                 local_init_done_from_the_frame_buffer,
                 local_refresh_ack_from_the_frame_buffer,
                 local_wdata_req_from_the_frame_buffer,
                 mem_addr_from_the_frame_buffer,
                 mem_ba_from_the_frame_buffer,
                 mem_cas_n_from_the_frame_buffer,
                 mem_cke_from_the_frame_buffer,
                 mem_clk_n_to_and_from_the_frame_buffer,
                 mem_clk_to_and_from_the_frame_buffer,
                 mem_cs_n_from_the_frame_buffer,
                 mem_dm_from_the_frame_buffer,
                 mem_dq_to_and_from_the_frame_buffer,
                 mem_dqs_to_and_from_the_frame_buffer,
                 mem_ras_n_from_the_frame_buffer,
                 mem_we_n_from_the_frame_buffer,
                 reset_phy_clk_n_from_the_frame_buffer,

                // the_lcd_i2c_cs
                 out_port_from_the_lcd_i2c_cs,

                // the_lcd_i2c_dat
                 bidir_port_to_and_from_the_lcd_i2c_dat,

                // the_lcd_i2c_scl
                 out_port_from_the_lcd_i2c_scl,

                // the_lcd_video_sequencer
                 DEN_from_the_lcd_video_sequencer,
                 HD_from_the_lcd_video_sequencer,
                 RGB_OUT_from_the_lcd_video_sequencer,
                 VD_from_the_lcd_video_sequencer,

                // the_pio_id_eeprom_dat
                 bidir_port_to_and_from_the_pio_id_eeprom_dat,

                // the_pio_id_eeprom_scl
                 out_port_from_the_pio_id_eeprom_scl,

                // the_push_buttons
                 in_port_to_the_push_buttons,

                // the_touchPanel_irq_n
                 in_port_to_the_touchPanel_irq_n,

                // the_touchPanel_spi
                 MISO_to_the_touchPanel_spi,
                 MOSI_from_the_touchPanel_spi,
                 SCLK_from_the_touchPanel_spi,
                 SS_n_from_the_touchPanel_spi,

                // the_tristate_bridge_avalon_slave
                 adsc_n_to_the_ssram,
                 bw_n_to_the_ssram,
                 bwe_n_to_the_ssram,
                 chipenable1_n_to_the_ssram,
                 outputenable_n_to_the_ssram,
                 read_n_to_the_flash,
                 reset_n_to_the_ssram,
                 select_n_to_the_flash,
                 tristate_bridge_address,
                 tristate_bridge_data,
                 write_n_to_the_flash
              )
;

  output           DEN_from_the_lcd_video_sequencer;
  output           HD_from_the_lcd_video_sequencer;
  output           MOSI_from_the_touchPanel_spi;
  output  [  7: 0] RGB_OUT_from_the_lcd_video_sequencer;
  output           SCLK_from_the_touchPanel_spi;
  output           SS_n_from_the_touchPanel_spi;
  output           VD_from_the_lcd_video_sequencer;
  output           adsc_n_to_the_ssram;
  inout            bidir_port_to_and_from_the_lcd_i2c_dat;
  inout            bidir_port_to_and_from_the_pio_id_eeprom_dat;
  output  [  3: 0] bw_n_to_the_ssram;
  output           bwe_n_to_the_ssram;
  output           chipenable1_n_to_the_ssram;
  output           frame_buffer_aux_full_rate_clk_out;
  output           frame_buffer_aux_half_rate_clk_out;
  output           frame_buffer_phy_clk_out;
  output           local_init_done_from_the_frame_buffer;
  output           local_refresh_ack_from_the_frame_buffer;
  output           local_wdata_req_from_the_frame_buffer;
  output  [ 12: 0] mem_addr_from_the_frame_buffer;
  output  [  1: 0] mem_ba_from_the_frame_buffer;
  output           mem_cas_n_from_the_frame_buffer;
  output           mem_cke_from_the_frame_buffer;
  inout            mem_clk_n_to_and_from_the_frame_buffer;
  inout            mem_clk_to_and_from_the_frame_buffer;
  output           mem_cs_n_from_the_frame_buffer;
  output  [  1: 0] mem_dm_from_the_frame_buffer;
  inout   [ 15: 0] mem_dq_to_and_from_the_frame_buffer;
  inout   [  1: 0] mem_dqs_to_and_from_the_frame_buffer;
  output           mem_ras_n_from_the_frame_buffer;
  output           mem_we_n_from_the_frame_buffer;
  output           out_port_from_the_lcd_i2c_cs;
  output           out_port_from_the_lcd_i2c_scl;
  output           out_port_from_the_pio_id_eeprom_scl;
  output           outputenable_n_to_the_ssram;
  output           read_n_to_the_flash;
  output           reset_n_to_the_ssram;
  output           reset_phy_clk_n_from_the_frame_buffer;
  output           select_n_to_the_flash;
  output  [ 23: 0] tristate_bridge_address;
  inout   [ 31: 0] tristate_bridge_data;
  output           write_n_to_the_flash;
  input            MISO_to_the_touchPanel_spi;
  input            ext_clk_one;
  input            global_reset_n_to_the_frame_buffer;
  input   [  3: 0] in_port_to_the_push_buttons;
  input            in_port_to_the_touchPanel_irq_n;
  input            reset_n;
  input            slow_clk;
  input            system_clk;
  input            video_clk;

  wire             DEN_from_the_lcd_video_sequencer;
  wire             HD_from_the_lcd_video_sequencer;
  wire             MOSI_from_the_touchPanel_spi;
  wire    [  7: 0] RGB_OUT_from_the_lcd_video_sequencer;
  wire             SCLK_from_the_touchPanel_spi;
  wire             SS_n_from_the_touchPanel_spi;
  wire             VD_from_the_lcd_video_sequencer;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave;
  wire    [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata;
  wire    [  3: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n;
  wire             accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa;
  wire             adsc_n_to_the_ssram;
  wire             bidir_port_to_and_from_the_lcd_i2c_dat;
  wire             bidir_port_to_and_from_the_pio_id_eeprom_dat;
  wire    [  3: 0] bw_n_to_the_ssram;
  wire             bwe_n_to_the_ssram;
  wire             chipenable1_n_to_the_ssram;
  wire    [ 10: 0] clock_crossing_bridge_m1_address;
  wire    [ 10: 0] clock_crossing_bridge_m1_address_to_slave;
  wire    [  3: 0] clock_crossing_bridge_m1_byteenable;
  wire             clock_crossing_bridge_m1_endofpacket;
  wire             clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_granted_push_buttons_s1;
  wire             clock_crossing_bridge_m1_granted_sysid_control_slave;
  wire             clock_crossing_bridge_m1_granted_system_tick_s1;
  wire             clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_latency_counter;
  wire    [  8: 0] clock_crossing_bridge_m1_nativeaddress;
  wire             clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_qualified_request_push_buttons_s1;
  wire             clock_crossing_bridge_m1_qualified_request_sysid_control_slave;
  wire             clock_crossing_bridge_m1_qualified_request_system_tick_s1;
  wire             clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_read;
  wire             clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_push_buttons_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_sysid_control_slave;
  wire             clock_crossing_bridge_m1_read_data_valid_system_tick_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port;
  wire    [ 31: 0] clock_crossing_bridge_m1_readdata;
  wire             clock_crossing_bridge_m1_readdatavalid;
  wire             clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1;
  wire             clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1;
  wire             clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1;
  wire             clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1;
  wire             clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1;
  wire             clock_crossing_bridge_m1_requests_push_buttons_s1;
  wire             clock_crossing_bridge_m1_requests_sysid_control_slave;
  wire             clock_crossing_bridge_m1_requests_system_tick_s1;
  wire             clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1;
  wire             clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port;
  wire             clock_crossing_bridge_m1_reset_n;
  wire             clock_crossing_bridge_m1_waitrequest;
  wire             clock_crossing_bridge_m1_write;
  wire    [ 31: 0] clock_crossing_bridge_m1_writedata;
  wire    [  8: 0] clock_crossing_bridge_s1_address;
  wire    [  3: 0] clock_crossing_bridge_s1_byteenable;
  wire             clock_crossing_bridge_s1_endofpacket;
  wire             clock_crossing_bridge_s1_endofpacket_from_sa;
  wire    [  8: 0] clock_crossing_bridge_s1_nativeaddress;
  wire             clock_crossing_bridge_s1_read;
  wire    [ 31: 0] clock_crossing_bridge_s1_readdata;
  wire    [ 31: 0] clock_crossing_bridge_s1_readdata_from_sa;
  wire             clock_crossing_bridge_s1_readdatavalid;
  wire             clock_crossing_bridge_s1_reset_n;
  wire             clock_crossing_bridge_s1_waitrequest;
  wire             clock_crossing_bridge_s1_waitrequest_from_sa;
  wire             clock_crossing_bridge_s1_write;
  wire    [ 31: 0] clock_crossing_bridge_s1_writedata;
  wire    [  7: 0] colour_lookup_table_s1_address;
  wire    [  3: 0] colour_lookup_table_s1_byteenable;
  wire             colour_lookup_table_s1_chipselect;
  wire             colour_lookup_table_s1_clken;
  wire    [ 31: 0] colour_lookup_table_s1_readdata;
  wire    [ 31: 0] colour_lookup_table_s1_readdata_from_sa;
  wire             colour_lookup_table_s1_reset;
  wire             colour_lookup_table_s1_write;
  wire    [ 31: 0] colour_lookup_table_s1_writedata;
  wire    [  7: 0] colour_lookup_table_s2_address;
  wire    [  3: 0] colour_lookup_table_s2_byteenable;
  wire             colour_lookup_table_s2_chipselect;
  wire             colour_lookup_table_s2_clken;
  wire    [ 31: 0] colour_lookup_table_s2_readdata;
  wire    [ 31: 0] colour_lookup_table_s2_readdata_from_sa;
  wire             colour_lookup_table_s2_reset;
  wire             colour_lookup_table_s2_write;
  wire    [ 31: 0] colour_lookup_table_s2_writedata;
  wire    [ 27: 0] cpu_data_master_address;
  wire    [ 27: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_granted_pipeline_bridge_s1;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_latency_counter;
  wire             cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_qualified_request_pipeline_bridge_s1;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0;
  wire             cpu_data_master_requests_pipeline_bridge_s1;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 26: 0] cpu_instruction_master_address;
  wire    [ 26: 0] cpu_instruction_master_address_to_slave;
  wire             cpu_instruction_master_granted_pipeline_bridge_s1;
  wire             cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_pipeline_bridge_s1;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_pipeline_bridge_s1;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire             d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer;
  wire             d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer;
  wire             d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer;
  wire             d1_clock_crossing_bridge_s1_end_xfer;
  wire             d1_colour_lookup_table_s1_end_xfer;
  wire             d1_colour_lookup_table_s2_end_xfer;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer;
  wire             d1_descriptor_memory_s1_end_xfer;
  wire             d1_descriptor_memory_s2_end_xfer;
  wire             d1_flash_ssram_pipeline_bridge_s1_end_xfer;
  wire             d1_frame_buffer_pipeline_bridge_s1_end_xfer;
  wire             d1_frame_buffer_s1_end_xfer;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_lcd_i2c_cs_s1_end_xfer;
  wire             d1_lcd_i2c_dat_s1_end_xfer;
  wire             d1_lcd_i2c_scl_s1_end_xfer;
  wire             d1_lcd_sgdma_csr_end_xfer;
  wire             d1_pio_id_eeprom_dat_s1_end_xfer;
  wire             d1_pio_id_eeprom_scl_s1_end_xfer;
  wire             d1_pipeline_bridge_s1_end_xfer;
  wire             d1_push_buttons_s1_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             d1_system_tick_s1_end_xfer;
  wire             d1_touchPanel_irq_n_s1_end_xfer;
  wire             d1_touchPanel_spi_spi_control_port_end_xfer;
  wire             d1_tristate_bridge_avalon_slave_end_xfer;
  wire    [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address;
  wire    [ 24: 0] ddr_sdram_clock_crossing_bridge_m1_address_to_slave;
  wire    [  3: 0] ddr_sdram_clock_crossing_bridge_m1_byteenable;
  wire             ddr_sdram_clock_crossing_bridge_m1_endofpacket;
  wire             ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_latency_counter;
  wire    [ 22: 0] ddr_sdram_clock_crossing_bridge_m1_nativeaddress;
  wire             ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_read;
  wire             ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_readdata;
  wire             ddr_sdram_clock_crossing_bridge_m1_readdatavalid;
  wire             ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1;
  wire             ddr_sdram_clock_crossing_bridge_m1_reset_n;
  wire             ddr_sdram_clock_crossing_bridge_m1_waitrequest;
  wire             ddr_sdram_clock_crossing_bridge_m1_write;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_m1_writedata;
  wire    [ 22: 0] ddr_sdram_clock_crossing_bridge_s1_address;
  wire    [  3: 0] ddr_sdram_clock_crossing_bridge_s1_byteenable;
  wire             ddr_sdram_clock_crossing_bridge_s1_endofpacket;
  wire             ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa;
  wire    [ 22: 0] ddr_sdram_clock_crossing_bridge_s1_nativeaddress;
  wire             ddr_sdram_clock_crossing_bridge_s1_read;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_readdata;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa;
  wire             ddr_sdram_clock_crossing_bridge_s1_readdatavalid;
  wire             ddr_sdram_clock_crossing_bridge_s1_reset_n;
  wire             ddr_sdram_clock_crossing_bridge_s1_waitrequest;
  wire             ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa;
  wire             ddr_sdram_clock_crossing_bridge_s1_write;
  wire    [ 31: 0] ddr_sdram_clock_crossing_bridge_s1_writedata;
  wire    [  9: 0] descriptor_memory_s1_address;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire             descriptor_memory_s1_clken;
  wire    [ 31: 0] descriptor_memory_s1_readdata;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  wire             descriptor_memory_s1_reset;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  wire    [  9: 0] descriptor_memory_s2_address;
  wire    [  3: 0] descriptor_memory_s2_byteenable;
  wire             descriptor_memory_s2_chipselect;
  wire             descriptor_memory_s2_clken;
  wire    [ 31: 0] descriptor_memory_s2_readdata;
  wire    [ 31: 0] descriptor_memory_s2_readdata_from_sa;
  wire             descriptor_memory_s2_reset;
  wire             descriptor_memory_s2_write;
  wire    [ 31: 0] descriptor_memory_s2_writedata;
  wire             dummy_master_inst_granted_colour_lookup_table_s2;
  wire    [ 31: 0] dummy_master_inst_m0_address;
  wire    [ 31: 0] dummy_master_inst_m0_address_to_slave;
  wire             dummy_master_inst_m0_waitrequest;
  wire             dummy_master_inst_m0_write;
  wire    [ 31: 0] dummy_master_inst_m0_writedata;
  wire             dummy_master_inst_qualified_request_colour_lookup_table_s2;
  wire             dummy_master_inst_requests_colour_lookup_table_s2;
  wire             ext_clk_one_reset_n;
  wire             flash_s1_wait_counter_eq_0;
  wire    [ 24: 0] flash_ssram_pipeline_bridge_m1_address;
  wire    [ 24: 0] flash_ssram_pipeline_bridge_m1_address_to_slave;
  wire             flash_ssram_pipeline_bridge_m1_burstcount;
  wire    [ 31: 0] flash_ssram_pipeline_bridge_m1_byteenable;
  wire    [  1: 0] flash_ssram_pipeline_bridge_m1_byteenable_flash_s1;
  wire    [  3: 0] flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1;
  wire             flash_ssram_pipeline_bridge_m1_chipselect;
  wire    [  4: 0] flash_ssram_pipeline_bridge_m1_dbs_address;
  wire    [ 15: 0] flash_ssram_pipeline_bridge_m1_dbs_write_16;
  wire    [ 31: 0] flash_ssram_pipeline_bridge_m1_dbs_write_32;
  wire             flash_ssram_pipeline_bridge_m1_debugaccess;
  wire             flash_ssram_pipeline_bridge_m1_endofpacket;
  wire             flash_ssram_pipeline_bridge_m1_granted_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_granted_ssram_s1;
  wire    [  2: 0] flash_ssram_pipeline_bridge_m1_latency_counter;
  wire             flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1;
  wire             flash_ssram_pipeline_bridge_m1_read;
  wire             flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1;
  wire    [255: 0] flash_ssram_pipeline_bridge_m1_readdata;
  wire             flash_ssram_pipeline_bridge_m1_readdatavalid;
  wire             flash_ssram_pipeline_bridge_m1_requests_flash_s1;
  wire             flash_ssram_pipeline_bridge_m1_requests_ssram_s1;
  wire             flash_ssram_pipeline_bridge_m1_waitrequest;
  wire             flash_ssram_pipeline_bridge_m1_write;
  wire    [255: 0] flash_ssram_pipeline_bridge_m1_writedata;
  wire    [ 19: 0] flash_ssram_pipeline_bridge_s1_address;
  wire             flash_ssram_pipeline_bridge_s1_arbiterlock;
  wire             flash_ssram_pipeline_bridge_s1_arbiterlock2;
  wire             flash_ssram_pipeline_bridge_s1_burstcount;
  wire    [ 31: 0] flash_ssram_pipeline_bridge_s1_byteenable;
  wire             flash_ssram_pipeline_bridge_s1_chipselect;
  wire             flash_ssram_pipeline_bridge_s1_debugaccess;
  wire             flash_ssram_pipeline_bridge_s1_endofpacket;
  wire             flash_ssram_pipeline_bridge_s1_endofpacket_from_sa;
  wire    [ 19: 0] flash_ssram_pipeline_bridge_s1_nativeaddress;
  wire             flash_ssram_pipeline_bridge_s1_read;
  wire    [255: 0] flash_ssram_pipeline_bridge_s1_readdata;
  wire    [255: 0] flash_ssram_pipeline_bridge_s1_readdata_from_sa;
  wire             flash_ssram_pipeline_bridge_s1_readdatavalid;
  wire             flash_ssram_pipeline_bridge_s1_reset_n;
  wire             flash_ssram_pipeline_bridge_s1_waitrequest;
  wire             flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
  wire             flash_ssram_pipeline_bridge_s1_write;
  wire    [255: 0] flash_ssram_pipeline_bridge_s1_writedata;
  wire             frame_buffer_aux_full_rate_clk_out;
  wire             frame_buffer_aux_half_rate_clk_out;
  wire             frame_buffer_phy_clk_out;
  wire             frame_buffer_phy_clk_out_reset_n;
  wire    [ 24: 0] frame_buffer_pipeline_bridge_m1_address;
  wire    [ 24: 0] frame_buffer_pipeline_bridge_m1_address_to_slave;
  wire             frame_buffer_pipeline_bridge_m1_burstcount;
  wire    [  3: 0] frame_buffer_pipeline_bridge_m1_byteenable;
  wire             frame_buffer_pipeline_bridge_m1_chipselect;
  wire             frame_buffer_pipeline_bridge_m1_debugaccess;
  wire             frame_buffer_pipeline_bridge_m1_endofpacket;
  wire             frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_latency_counter;
  wire             frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_read;
  wire             frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_m1_readdata;
  wire             frame_buffer_pipeline_bridge_m1_readdatavalid;
  wire             frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1;
  wire             frame_buffer_pipeline_bridge_m1_waitrequest;
  wire             frame_buffer_pipeline_bridge_m1_write;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_m1_writedata;
  wire    [ 22: 0] frame_buffer_pipeline_bridge_s1_address;
  wire             frame_buffer_pipeline_bridge_s1_arbiterlock;
  wire             frame_buffer_pipeline_bridge_s1_arbiterlock2;
  wire             frame_buffer_pipeline_bridge_s1_burstcount;
  wire    [  3: 0] frame_buffer_pipeline_bridge_s1_byteenable;
  wire             frame_buffer_pipeline_bridge_s1_chipselect;
  wire             frame_buffer_pipeline_bridge_s1_debugaccess;
  wire             frame_buffer_pipeline_bridge_s1_endofpacket;
  wire             frame_buffer_pipeline_bridge_s1_endofpacket_from_sa;
  wire    [ 22: 0] frame_buffer_pipeline_bridge_s1_nativeaddress;
  wire             frame_buffer_pipeline_bridge_s1_read;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_s1_readdata_from_sa;
  wire             frame_buffer_pipeline_bridge_s1_readdatavalid;
  wire             frame_buffer_pipeline_bridge_s1_reset_n;
  wire             frame_buffer_pipeline_bridge_s1_waitrequest;
  wire             frame_buffer_pipeline_bridge_s1_waitrequest_from_sa;
  wire             frame_buffer_pipeline_bridge_s1_write;
  wire    [ 31: 0] frame_buffer_pipeline_bridge_s1_writedata;
  wire    [ 22: 0] frame_buffer_s1_address;
  wire             frame_buffer_s1_beginbursttransfer;
  wire    [  1: 0] frame_buffer_s1_burstcount;
  wire    [  3: 0] frame_buffer_s1_byteenable;
  wire             frame_buffer_s1_read;
  wire    [ 31: 0] frame_buffer_s1_readdata;
  wire    [ 31: 0] frame_buffer_s1_readdata_from_sa;
  wire             frame_buffer_s1_readdatavalid;
  wire             frame_buffer_s1_resetrequest_n;
  wire             frame_buffer_s1_resetrequest_n_from_sa;
  wire             frame_buffer_s1_waitrequest_n;
  wire             frame_buffer_s1_waitrequest_n_from_sa;
  wire             frame_buffer_s1_write;
  wire    [ 31: 0] frame_buffer_s1_writedata;
  wire    [ 31: 0] incoming_tristate_bridge_data;
  wire    [ 15: 0] incoming_tristate_bridge_data_with_Xs_converted_to_0;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire    [  7: 0] lcd_data_format_adapter_1_in_data;
  wire             lcd_data_format_adapter_1_in_endofpacket;
  wire             lcd_data_format_adapter_1_in_ready;
  wire             lcd_data_format_adapter_1_in_ready_from_sa;
  wire             lcd_data_format_adapter_1_in_reset_n;
  wire             lcd_data_format_adapter_1_in_startofpacket;
  wire             lcd_data_format_adapter_1_in_valid;
  wire    [  7: 0] lcd_data_format_adapter_1_out_data;
  wire             lcd_data_format_adapter_1_out_empty;
  wire             lcd_data_format_adapter_1_out_endofpacket;
  wire             lcd_data_format_adapter_1_out_ready;
  wire             lcd_data_format_adapter_1_out_startofpacket;
  wire             lcd_data_format_adapter_1_out_valid;
  wire    [ 23: 0] lcd_data_format_adapter_in_data;
  wire    [  1: 0] lcd_data_format_adapter_in_empty;
  wire             lcd_data_format_adapter_in_endofpacket;
  wire             lcd_data_format_adapter_in_ready;
  wire             lcd_data_format_adapter_in_ready_from_sa;
  wire             lcd_data_format_adapter_in_reset_n;
  wire             lcd_data_format_adapter_in_startofpacket;
  wire             lcd_data_format_adapter_in_valid;
  wire    [  7: 0] lcd_data_format_adapter_out_data;
  wire             lcd_data_format_adapter_out_endofpacket;
  wire             lcd_data_format_adapter_out_ready;
  wire             lcd_data_format_adapter_out_startofpacket;
  wire             lcd_data_format_adapter_out_valid;
  wire    [  1: 0] lcd_i2c_cs_s1_address;
  wire             lcd_i2c_cs_s1_chipselect;
  wire    [ 31: 0] lcd_i2c_cs_s1_readdata;
  wire    [ 31: 0] lcd_i2c_cs_s1_readdata_from_sa;
  wire             lcd_i2c_cs_s1_reset_n;
  wire             lcd_i2c_cs_s1_write_n;
  wire    [ 31: 0] lcd_i2c_cs_s1_writedata;
  wire    [  1: 0] lcd_i2c_dat_s1_address;
  wire             lcd_i2c_dat_s1_chipselect;
  wire    [ 31: 0] lcd_i2c_dat_s1_readdata;
  wire    [ 31: 0] lcd_i2c_dat_s1_readdata_from_sa;
  wire             lcd_i2c_dat_s1_reset_n;
  wire             lcd_i2c_dat_s1_write_n;
  wire    [ 31: 0] lcd_i2c_dat_s1_writedata;
  wire    [  1: 0] lcd_i2c_scl_s1_address;
  wire             lcd_i2c_scl_s1_chipselect;
  wire    [ 31: 0] lcd_i2c_scl_s1_readdata;
  wire    [ 31: 0] lcd_i2c_scl_s1_readdata_from_sa;
  wire             lcd_i2c_scl_s1_reset_n;
  wire             lcd_i2c_scl_s1_write_n;
  wire    [ 31: 0] lcd_i2c_scl_s1_writedata;
  wire    [  7: 0] lcd_on_chip_memory_fifo_in_data;
  wire             lcd_on_chip_memory_fifo_in_endofpacket;
  wire             lcd_on_chip_memory_fifo_in_ready;
  wire             lcd_on_chip_memory_fifo_in_ready_from_sa;
  wire             lcd_on_chip_memory_fifo_in_reset_n;
  wire             lcd_on_chip_memory_fifo_in_startofpacket;
  wire             lcd_on_chip_memory_fifo_in_valid;
  wire    [  7: 0] lcd_on_chip_memory_fifo_out_data;
  wire             lcd_on_chip_memory_fifo_out_endofpacket;
  wire             lcd_on_chip_memory_fifo_out_ready;
  wire             lcd_on_chip_memory_fifo_out_reset_n;
  wire             lcd_on_chip_memory_fifo_out_startofpacket;
  wire             lcd_on_chip_memory_fifo_out_valid;
  wire    [ 31: 0] lcd_pixel_converter_in_data;
  wire    [  1: 0] lcd_pixel_converter_in_empty;
  wire             lcd_pixel_converter_in_endofpacket;
  wire             lcd_pixel_converter_in_ready;
  wire             lcd_pixel_converter_in_ready_from_sa;
  wire             lcd_pixel_converter_in_reset_n;
  wire             lcd_pixel_converter_in_startofpacket;
  wire             lcd_pixel_converter_in_valid;
  wire    [ 23: 0] lcd_pixel_converter_out_data;
  wire    [  1: 0] lcd_pixel_converter_out_empty;
  wire             lcd_pixel_converter_out_endofpacket;
  wire             lcd_pixel_converter_out_ready;
  wire             lcd_pixel_converter_out_startofpacket;
  wire             lcd_pixel_converter_out_valid;
  wire    [  3: 0] lcd_sgdma_csr_address;
  wire             lcd_sgdma_csr_chipselect;
  wire             lcd_sgdma_csr_irq;
  wire             lcd_sgdma_csr_irq_from_sa;
  wire             lcd_sgdma_csr_read;
  wire    [ 31: 0] lcd_sgdma_csr_readdata;
  wire    [ 31: 0] lcd_sgdma_csr_readdata_from_sa;
  wire             lcd_sgdma_csr_reset_n;
  wire             lcd_sgdma_csr_write;
  wire    [ 31: 0] lcd_sgdma_csr_writedata;
  wire    [ 31: 0] lcd_sgdma_descriptor_read_address;
  wire    [ 31: 0] lcd_sgdma_descriptor_read_address_to_slave;
  wire             lcd_sgdma_descriptor_read_granted_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_latency_counter;
  wire             lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_read;
  wire             lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2;
  wire    [ 31: 0] lcd_sgdma_descriptor_read_readdata;
  wire             lcd_sgdma_descriptor_read_readdatavalid;
  wire             lcd_sgdma_descriptor_read_requests_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_read_waitrequest;
  wire    [ 31: 0] lcd_sgdma_descriptor_write_address;
  wire    [ 31: 0] lcd_sgdma_descriptor_write_address_to_slave;
  wire             lcd_sgdma_descriptor_write_granted_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_requests_descriptor_memory_s2;
  wire             lcd_sgdma_descriptor_write_waitrequest;
  wire             lcd_sgdma_descriptor_write_write;
  wire    [ 31: 0] lcd_sgdma_descriptor_write_writedata;
  wire    [ 31: 0] lcd_sgdma_m_read_address;
  wire    [ 31: 0] lcd_sgdma_m_read_address_to_slave;
  wire             lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_latency_counter;
  wire             lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_read;
  wire             lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  wire    [ 31: 0] lcd_sgdma_m_read_readdata;
  wire             lcd_sgdma_m_read_readdatavalid;
  wire             lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1;
  wire             lcd_sgdma_m_read_waitrequest;
  wire    [ 31: 0] lcd_sgdma_out_data;
  wire    [  1: 0] lcd_sgdma_out_empty;
  wire             lcd_sgdma_out_endofpacket;
  wire             lcd_sgdma_out_ready;
  wire             lcd_sgdma_out_startofpacket;
  wire             lcd_sgdma_out_valid;
  wire    [  7: 0] lcd_ta_fifo_to_sequencer_in_data;
  wire             lcd_ta_fifo_to_sequencer_in_endofpacket;
  wire             lcd_ta_fifo_to_sequencer_in_ready;
  wire             lcd_ta_fifo_to_sequencer_in_ready_from_sa;
  wire             lcd_ta_fifo_to_sequencer_in_reset_n;
  wire             lcd_ta_fifo_to_sequencer_in_startofpacket;
  wire             lcd_ta_fifo_to_sequencer_in_valid;
  wire    [  7: 0] lcd_ta_fifo_to_sequencer_out_data;
  wire             lcd_ta_fifo_to_sequencer_out_endofpacket;
  wire             lcd_ta_fifo_to_sequencer_out_ready;
  wire             lcd_ta_fifo_to_sequencer_out_startofpacket;
  wire             lcd_ta_fifo_to_sequencer_out_valid;
  wire    [  7: 0] lcd_ta_formatter_to_fifo_in_data;
  wire             lcd_ta_formatter_to_fifo_in_endofpacket;
  wire             lcd_ta_formatter_to_fifo_in_ready;
  wire             lcd_ta_formatter_to_fifo_in_ready_from_sa;
  wire             lcd_ta_formatter_to_fifo_in_reset_n;
  wire             lcd_ta_formatter_to_fifo_in_startofpacket;
  wire             lcd_ta_formatter_to_fifo_in_valid;
  wire    [  7: 0] lcd_ta_formatter_to_fifo_out_data;
  wire             lcd_ta_formatter_to_fifo_out_endofpacket;
  wire             lcd_ta_formatter_to_fifo_out_ready;
  wire             lcd_ta_formatter_to_fifo_out_startofpacket;
  wire             lcd_ta_formatter_to_fifo_out_valid;
  wire    [  7: 0] lcd_video_sequencer_in_data;
  wire             lcd_video_sequencer_in_empty;
  wire             lcd_video_sequencer_in_endofpacket;
  wire             lcd_video_sequencer_in_ready;
  wire             lcd_video_sequencer_in_ready_from_sa;
  wire             lcd_video_sequencer_in_reset_n;
  wire             lcd_video_sequencer_in_startofpacket;
  wire             lcd_video_sequencer_in_valid;
  wire             local_init_done_from_the_frame_buffer;
  wire             local_refresh_ack_from_the_frame_buffer;
  wire             local_wdata_req_from_the_frame_buffer;
  wire    [ 12: 0] mem_addr_from_the_frame_buffer;
  wire    [  1: 0] mem_ba_from_the_frame_buffer;
  wire             mem_cas_n_from_the_frame_buffer;
  wire             mem_cke_from_the_frame_buffer;
  wire             mem_clk_n_to_and_from_the_frame_buffer;
  wire             mem_clk_to_and_from_the_frame_buffer;
  wire             mem_cs_n_from_the_frame_buffer;
  wire    [  1: 0] mem_dm_from_the_frame_buffer;
  wire    [ 15: 0] mem_dq_to_and_from_the_frame_buffer;
  wire    [  1: 0] mem_dqs_to_and_from_the_frame_buffer;
  wire             mem_ras_n_from_the_frame_buffer;
  wire             mem_we_n_from_the_frame_buffer;
  wire             out_clk_frame_buffer_aux_full_rate_clk;
  wire             out_clk_frame_buffer_aux_half_rate_clk;
  wire             out_clk_frame_buffer_phy_clk;
  wire             out_port_from_the_lcd_i2c_cs;
  wire             out_port_from_the_lcd_i2c_scl;
  wire             out_port_from_the_pio_id_eeprom_scl;
  wire             outputenable_n_to_the_ssram;
  wire    [  1: 0] pio_id_eeprom_dat_s1_address;
  wire             pio_id_eeprom_dat_s1_chipselect;
  wire    [ 31: 0] pio_id_eeprom_dat_s1_readdata;
  wire    [ 31: 0] pio_id_eeprom_dat_s1_readdata_from_sa;
  wire             pio_id_eeprom_dat_s1_reset_n;
  wire             pio_id_eeprom_dat_s1_write_n;
  wire    [ 31: 0] pio_id_eeprom_dat_s1_writedata;
  wire    [  1: 0] pio_id_eeprom_scl_s1_address;
  wire             pio_id_eeprom_scl_s1_chipselect;
  wire    [ 31: 0] pio_id_eeprom_scl_s1_readdata;
  wire    [ 31: 0] pio_id_eeprom_scl_s1_readdata_from_sa;
  wire             pio_id_eeprom_scl_s1_reset_n;
  wire             pio_id_eeprom_scl_s1_write_n;
  wire    [ 31: 0] pio_id_eeprom_scl_s1_writedata;
  wire    [ 26: 0] pipeline_bridge_m1_address;
  wire    [ 26: 0] pipeline_bridge_m1_address_to_slave;
  wire             pipeline_bridge_m1_burstcount;
  wire    [  3: 0] pipeline_bridge_m1_byteenable;
  wire             pipeline_bridge_m1_chipselect;
  wire             pipeline_bridge_m1_debugaccess;
  wire             pipeline_bridge_m1_endofpacket;
  wire             pipeline_bridge_m1_granted_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_granted_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_granted_descriptor_memory_s1;
  wire             pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_granted_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_latency_counter;
  wire             pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_qualified_request_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_qualified_request_descriptor_memory_s1;
  wire             pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_qualified_request_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_read;
  wire             pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register;
  wire             pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_read_data_valid_descriptor_memory_s1;
  wire             pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  wire             pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register;
  wire             pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr;
  wire    [ 31: 0] pipeline_bridge_m1_readdata;
  wire             pipeline_bridge_m1_readdatavalid;
  wire             pipeline_bridge_m1_requests_clock_crossing_bridge_s1;
  wire             pipeline_bridge_m1_requests_colour_lookup_table_s1;
  wire             pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_requests_descriptor_memory_s1;
  wire             pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1;
  wire             pipeline_bridge_m1_requests_lcd_sgdma_csr;
  wire             pipeline_bridge_m1_waitrequest;
  wire             pipeline_bridge_m1_write;
  wire    [ 31: 0] pipeline_bridge_m1_writedata;
  wire    [ 24: 0] pipeline_bridge_s1_address;
  wire             pipeline_bridge_s1_arbiterlock;
  wire             pipeline_bridge_s1_arbiterlock2;
  wire             pipeline_bridge_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_s1_byteenable;
  wire             pipeline_bridge_s1_chipselect;
  wire             pipeline_bridge_s1_debugaccess;
  wire             pipeline_bridge_s1_endofpacket;
  wire             pipeline_bridge_s1_endofpacket_from_sa;
  wire    [ 24: 0] pipeline_bridge_s1_nativeaddress;
  wire             pipeline_bridge_s1_read;
  wire    [ 31: 0] pipeline_bridge_s1_readdata;
  wire    [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  wire             pipeline_bridge_s1_readdatavalid;
  wire             pipeline_bridge_s1_reset_n;
  wire             pipeline_bridge_s1_waitrequest;
  wire             pipeline_bridge_s1_waitrequest_from_sa;
  wire             pipeline_bridge_s1_write;
  wire    [ 31: 0] pipeline_bridge_s1_writedata;
  wire    [  1: 0] push_buttons_s1_address;
  wire             push_buttons_s1_chipselect;
  wire             push_buttons_s1_irq;
  wire             push_buttons_s1_irq_from_sa;
  wire    [ 31: 0] push_buttons_s1_readdata;
  wire    [ 31: 0] push_buttons_s1_readdata_from_sa;
  wire             push_buttons_s1_reset_n;
  wire             push_buttons_s1_write_n;
  wire    [ 31: 0] push_buttons_s1_writedata;
  wire             read_n_to_the_flash;
  wire             reset_n_sources;
  wire             reset_n_to_the_ssram;
  wire             reset_phy_clk_n_from_the_frame_buffer;
  wire             select_n_to_the_flash;
  wire             slow_clk_reset_n;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_clock;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             sysid_control_slave_reset_n;
  wire             system_clk_reset_n;
  wire    [  2: 0] system_tick_s1_address;
  wire             system_tick_s1_chipselect;
  wire             system_tick_s1_irq;
  wire             system_tick_s1_irq_from_sa;
  wire    [ 15: 0] system_tick_s1_readdata;
  wire    [ 15: 0] system_tick_s1_readdata_from_sa;
  wire             system_tick_s1_reset_n;
  wire             system_tick_s1_write_n;
  wire    [ 15: 0] system_tick_s1_writedata;
  wire    [  1: 0] touchPanel_irq_n_s1_address;
  wire             touchPanel_irq_n_s1_chipselect;
  wire             touchPanel_irq_n_s1_irq;
  wire             touchPanel_irq_n_s1_irq_from_sa;
  wire    [ 31: 0] touchPanel_irq_n_s1_readdata;
  wire    [ 31: 0] touchPanel_irq_n_s1_readdata_from_sa;
  wire             touchPanel_irq_n_s1_reset_n;
  wire             touchPanel_irq_n_s1_write_n;
  wire    [ 31: 0] touchPanel_irq_n_s1_writedata;
  wire    [  2: 0] touchPanel_spi_spi_control_port_address;
  wire             touchPanel_spi_spi_control_port_chipselect;
  wire             touchPanel_spi_spi_control_port_dataavailable;
  wire             touchPanel_spi_spi_control_port_dataavailable_from_sa;
  wire             touchPanel_spi_spi_control_port_endofpacket;
  wire             touchPanel_spi_spi_control_port_endofpacket_from_sa;
  wire             touchPanel_spi_spi_control_port_irq;
  wire             touchPanel_spi_spi_control_port_irq_from_sa;
  wire             touchPanel_spi_spi_control_port_read_n;
  wire    [ 15: 0] touchPanel_spi_spi_control_port_readdata;
  wire    [ 15: 0] touchPanel_spi_spi_control_port_readdata_from_sa;
  wire             touchPanel_spi_spi_control_port_readyfordata;
  wire             touchPanel_spi_spi_control_port_readyfordata_from_sa;
  wire             touchPanel_spi_spi_control_port_reset_n;
  wire             touchPanel_spi_spi_control_port_write_n;
  wire    [ 15: 0] touchPanel_spi_spi_control_port_writedata;
  wire    [ 23: 0] tristate_bridge_address;
  wire    [ 31: 0] tristate_bridge_data;
  wire             video_clk_reset_n;
  wire             write_n_to_the_flash;
  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address                           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq                               (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa                       (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n                           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata),
      .clk                                                                                                             (system_clk),
      .cpu_data_master_address_to_slave                                                                                (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0           (cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_latency_counter                                                                                 (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 (cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_read                                                                                            (cpu_data_master_read),
      .cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0   (cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register                                               (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register),
      .cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0          (cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_write                                                                                           (cpu_data_master_write),
      .cpu_data_master_writedata                                                                                       (cpu_data_master_writedata),
      .d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer                       (d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer),
      .reset_n                                                                                                         (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave                                                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write                                                                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address                                                                                       (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect                                                                                    (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata                                                                                      (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa                                                                              (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa),
      .clk                                                                                                                                                                      (system_clk),
      .d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer                                                                                   (d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer),
      .reset_n                                                                                                                                                                  (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave                                                                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read                                                                                                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer                                                                                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect                                                                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read                                                                                              (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata                                                                                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa                                                                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n                                                                                           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n                                                                                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa                                                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa),
      .clk                                                                                                                                                                                          (system_clk),
      .d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer                                                                                       (d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer),
      .reset_n                                                                                                                                                                                      (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush                                    (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported                 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read                                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata                                 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid                            (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n                            (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n),
      .clk                                                                                                                                                                    (system_clk),
      .colour_lookup_table_s2_readdata_from_sa                                                                                                                                (colour_lookup_table_s2_readdata_from_sa),
      .d1_colour_lookup_table_s2_end_xfer                                                                                                                                     (d1_colour_lookup_table_s2_end_xfer),
      .reset_n                                                                                                                                                                (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address                                           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n                                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata                                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata),
      .clk                                                                                                                                                                             (system_clk),
      .d1_frame_buffer_pipeline_bridge_s1_end_xfer                                                                                                                                     (d1_frame_buffer_pipeline_bridge_s1_end_xfer),
      .frame_buffer_pipeline_bridge_s1_waitrequest_from_sa                                                                                                                             (frame_buffer_pipeline_bridge_s1_waitrequest_from_sa),
      .reset_n                                                                                                                                                                         (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address                                                                                      (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave                                                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest                                                                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write                                                                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata                                                                                    (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata),
      .clk                                                                                                                                                                      (system_clk),
      .d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer                                                                                   (d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_end_xfer),
      .reset_n                                                                                                                                                                  (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_arbitrator the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address                                                                                                      (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave                                                                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read                                                                                                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata                                                                                                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n                                                                                                (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa                                                                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa                                                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n_from_sa),
      .clk                                                                                                                                                                                          (system_clk),
      .d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer                                                                                       (d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_end_xfer),
      .reset_n                                                                                                                                                                                      (system_clk_reset_n)
    );

  accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance the_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address0       (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush0         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read0          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata0      (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdata),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid0 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_readdatavalid),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n0 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_waitrequest_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address0       (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable0    (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n0 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_waitrequest_n),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write0         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata0     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata),
      .clk                                                                           (system_clk),
      .cpu_address0                                                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_address),
      .cpu_clk                                                                       (system_clk),
      .cpu_irq0                                                                      (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq),
      .cpu_readdata0                                                                 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_readdata),
      .cpu_readdata1                                                                 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata),
      .cpu_reset_n                                                                   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_reset_n),
      .cpu_select0                                                                   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_chipselect),
      .cpu_waitrequest_n0                                                            (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n),
      .cpu_write0                                                                    (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_write),
      .cpu_writedata0                                                                (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_writedata),
      .dummy_master_address                                                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_address),
      .dummy_master_waitrequest                                                      (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_waitrequest),
      .dummy_master_write                                                            (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_write),
      .dummy_master_writedata                                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_master_writedata),
      .dummy_slave_address                                                           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_address),
      .dummy_slave_chipselect                                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_chipselect),
      .dummy_slave_readdata                                                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata),
      .hw_draw_int_mandelbrot_begin0                                                 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_begintransfer),
      .hw_draw_int_mandelbrot_read0                                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_read),
      .hw_draw_int_mandelbrot_select0                                                (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_chipselect),
      .hw_draw_int_mandelbrot_waitrequest_n0                                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_waitrequest_n),
      .reset_n                                                                       (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_sub_hw_draw_int_mandelbrot0_reset_n),
      .slave_address0                                                                (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_address),
      .slave_read0                                                                   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_read),
      .slave_readdata0                                                               (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_readdata),
      .slave_waitrequest_n0                                                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_internal_master0_waitrequest_n)
    );

  clock_crossing_bridge_s1_arbitrator the_clock_crossing_bridge_s1
    (
      .clk                                                                               (system_clk),
      .clock_crossing_bridge_s1_address                                                  (clock_crossing_bridge_s1_address),
      .clock_crossing_bridge_s1_byteenable                                               (clock_crossing_bridge_s1_byteenable),
      .clock_crossing_bridge_s1_endofpacket                                              (clock_crossing_bridge_s1_endofpacket),
      .clock_crossing_bridge_s1_endofpacket_from_sa                                      (clock_crossing_bridge_s1_endofpacket_from_sa),
      .clock_crossing_bridge_s1_nativeaddress                                            (clock_crossing_bridge_s1_nativeaddress),
      .clock_crossing_bridge_s1_read                                                     (clock_crossing_bridge_s1_read),
      .clock_crossing_bridge_s1_readdata                                                 (clock_crossing_bridge_s1_readdata),
      .clock_crossing_bridge_s1_readdata_from_sa                                         (clock_crossing_bridge_s1_readdata_from_sa),
      .clock_crossing_bridge_s1_readdatavalid                                            (clock_crossing_bridge_s1_readdatavalid),
      .clock_crossing_bridge_s1_reset_n                                                  (clock_crossing_bridge_s1_reset_n),
      .clock_crossing_bridge_s1_waitrequest                                              (clock_crossing_bridge_s1_waitrequest),
      .clock_crossing_bridge_s1_waitrequest_from_sa                                      (clock_crossing_bridge_s1_waitrequest_from_sa),
      .clock_crossing_bridge_s1_write                                                    (clock_crossing_bridge_s1_write),
      .clock_crossing_bridge_s1_writedata                                                (clock_crossing_bridge_s1_writedata),
      .d1_clock_crossing_bridge_s1_end_xfer                                              (d1_clock_crossing_bridge_s1_end_xfer),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                     (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_clock_crossing_bridge_s1                               (pipeline_bridge_m1_granted_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1                     (pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1                       (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_requests_clock_crossing_bridge_s1                              (pipeline_bridge_m1_requests_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  clock_crossing_bridge_m1_arbitrator the_clock_crossing_bridge_m1
    (
      .clk                                                                        (slow_clk),
      .clock_crossing_bridge_m1_address                                           (clock_crossing_bridge_m1_address),
      .clock_crossing_bridge_m1_address_to_slave                                  (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_byteenable                                        (clock_crossing_bridge_m1_byteenable),
      .clock_crossing_bridge_m1_endofpacket                                       (clock_crossing_bridge_m1_endofpacket),
      .clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave               (clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1                             (clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1                            (clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1                            (clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1                      (clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1                      (clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_granted_push_buttons_s1                           (clock_crossing_bridge_m1_granted_push_buttons_s1),
      .clock_crossing_bridge_m1_granted_sysid_control_slave                       (clock_crossing_bridge_m1_granted_sysid_control_slave),
      .clock_crossing_bridge_m1_granted_system_tick_s1                            (clock_crossing_bridge_m1_granted_system_tick_s1),
      .clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1                       (clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port           (clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_latency_counter                                   (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave     (clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1                   (clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1                  (clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1                  (clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1            (clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1            (clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_qualified_request_push_buttons_s1                 (clock_crossing_bridge_m1_qualified_request_push_buttons_s1),
      .clock_crossing_bridge_m1_qualified_request_sysid_control_slave             (clock_crossing_bridge_m1_qualified_request_sysid_control_slave),
      .clock_crossing_bridge_m1_qualified_request_system_tick_s1                  (clock_crossing_bridge_m1_qualified_request_system_tick_s1),
      .clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1             (clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port (clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_read                                              (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave       (clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1                     (clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1                    (clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1                    (clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1              (clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1              (clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_read_data_valid_push_buttons_s1                   (clock_crossing_bridge_m1_read_data_valid_push_buttons_s1),
      .clock_crossing_bridge_m1_read_data_valid_sysid_control_slave               (clock_crossing_bridge_m1_read_data_valid_sysid_control_slave),
      .clock_crossing_bridge_m1_read_data_valid_system_tick_s1                    (clock_crossing_bridge_m1_read_data_valid_system_tick_s1),
      .clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1               (clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port   (clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_readdata                                          (clock_crossing_bridge_m1_readdata),
      .clock_crossing_bridge_m1_readdatavalid                                     (clock_crossing_bridge_m1_readdatavalid),
      .clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave              (clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1                            (clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1                           (clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1                           (clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1                     (clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1                     (clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_requests_push_buttons_s1                          (clock_crossing_bridge_m1_requests_push_buttons_s1),
      .clock_crossing_bridge_m1_requests_sysid_control_slave                      (clock_crossing_bridge_m1_requests_sysid_control_slave),
      .clock_crossing_bridge_m1_requests_system_tick_s1                           (clock_crossing_bridge_m1_requests_system_tick_s1),
      .clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1                      (clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port          (clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_reset_n                                           (clock_crossing_bridge_m1_reset_n),
      .clock_crossing_bridge_m1_waitrequest                                       (clock_crossing_bridge_m1_waitrequest),
      .clock_crossing_bridge_m1_write                                             (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                                         (clock_crossing_bridge_m1_writedata),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                    (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .d1_lcd_i2c_cs_s1_end_xfer                                                  (d1_lcd_i2c_cs_s1_end_xfer),
      .d1_lcd_i2c_dat_s1_end_xfer                                                 (d1_lcd_i2c_dat_s1_end_xfer),
      .d1_lcd_i2c_scl_s1_end_xfer                                                 (d1_lcd_i2c_scl_s1_end_xfer),
      .d1_pio_id_eeprom_dat_s1_end_xfer                                           (d1_pio_id_eeprom_dat_s1_end_xfer),
      .d1_pio_id_eeprom_scl_s1_end_xfer                                           (d1_pio_id_eeprom_scl_s1_end_xfer),
      .d1_push_buttons_s1_end_xfer                                                (d1_push_buttons_s1_end_xfer),
      .d1_sysid_control_slave_end_xfer                                            (d1_sysid_control_slave_end_xfer),
      .d1_system_tick_s1_end_xfer                                                 (d1_system_tick_s1_end_xfer),
      .d1_touchPanel_irq_n_s1_end_xfer                                            (d1_touchPanel_irq_n_s1_end_xfer),
      .d1_touchPanel_spi_spi_control_port_end_xfer                                (d1_touchPanel_spi_spi_control_port_end_xfer),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                               (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                            (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .lcd_i2c_cs_s1_readdata_from_sa                                             (lcd_i2c_cs_s1_readdata_from_sa),
      .lcd_i2c_dat_s1_readdata_from_sa                                            (lcd_i2c_dat_s1_readdata_from_sa),
      .lcd_i2c_scl_s1_readdata_from_sa                                            (lcd_i2c_scl_s1_readdata_from_sa),
      .pio_id_eeprom_dat_s1_readdata_from_sa                                      (pio_id_eeprom_dat_s1_readdata_from_sa),
      .pio_id_eeprom_scl_s1_readdata_from_sa                                      (pio_id_eeprom_scl_s1_readdata_from_sa),
      .push_buttons_s1_readdata_from_sa                                           (push_buttons_s1_readdata_from_sa),
      .reset_n                                                                    (slow_clk_reset_n),
      .sysid_control_slave_readdata_from_sa                                       (sysid_control_slave_readdata_from_sa),
      .system_tick_s1_readdata_from_sa                                            (system_tick_s1_readdata_from_sa),
      .touchPanel_irq_n_s1_readdata_from_sa                                       (touchPanel_irq_n_s1_readdata_from_sa),
      .touchPanel_spi_spi_control_port_endofpacket_from_sa                        (touchPanel_spi_spi_control_port_endofpacket_from_sa),
      .touchPanel_spi_spi_control_port_readdata_from_sa                           (touchPanel_spi_spi_control_port_readdata_from_sa)
    );

  clock_crossing_bridge the_clock_crossing_bridge
    (
      .master_address       (clock_crossing_bridge_m1_address),
      .master_byteenable    (clock_crossing_bridge_m1_byteenable),
      .master_clk           (slow_clk),
      .master_endofpacket   (clock_crossing_bridge_m1_endofpacket),
      .master_nativeaddress (clock_crossing_bridge_m1_nativeaddress),
      .master_read          (clock_crossing_bridge_m1_read),
      .master_readdata      (clock_crossing_bridge_m1_readdata),
      .master_readdatavalid (clock_crossing_bridge_m1_readdatavalid),
      .master_reset_n       (clock_crossing_bridge_m1_reset_n),
      .master_waitrequest   (clock_crossing_bridge_m1_waitrequest),
      .master_write         (clock_crossing_bridge_m1_write),
      .master_writedata     (clock_crossing_bridge_m1_writedata),
      .slave_address        (clock_crossing_bridge_s1_address),
      .slave_byteenable     (clock_crossing_bridge_s1_byteenable),
      .slave_clk            (system_clk),
      .slave_endofpacket    (clock_crossing_bridge_s1_endofpacket),
      .slave_nativeaddress  (clock_crossing_bridge_s1_nativeaddress),
      .slave_read           (clock_crossing_bridge_s1_read),
      .slave_readdata       (clock_crossing_bridge_s1_readdata),
      .slave_readdatavalid  (clock_crossing_bridge_s1_readdatavalid),
      .slave_reset_n        (clock_crossing_bridge_s1_reset_n),
      .slave_waitrequest    (clock_crossing_bridge_s1_waitrequest),
      .slave_write          (clock_crossing_bridge_s1_write),
      .slave_writedata      (clock_crossing_bridge_s1_writedata)
    );

  colour_lookup_table_s1_arbitrator the_colour_lookup_table_s1
    (
      .clk                                                                               (system_clk),
      .colour_lookup_table_s1_address                                                    (colour_lookup_table_s1_address),
      .colour_lookup_table_s1_byteenable                                                 (colour_lookup_table_s1_byteenable),
      .colour_lookup_table_s1_chipselect                                                 (colour_lookup_table_s1_chipselect),
      .colour_lookup_table_s1_clken                                                      (colour_lookup_table_s1_clken),
      .colour_lookup_table_s1_readdata                                                   (colour_lookup_table_s1_readdata),
      .colour_lookup_table_s1_readdata_from_sa                                           (colour_lookup_table_s1_readdata_from_sa),
      .colour_lookup_table_s1_reset                                                      (colour_lookup_table_s1_reset),
      .colour_lookup_table_s1_write                                                      (colour_lookup_table_s1_write),
      .colour_lookup_table_s1_writedata                                                  (colour_lookup_table_s1_writedata),
      .d1_colour_lookup_table_s1_end_xfer                                                (d1_colour_lookup_table_s1_end_xfer),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                     (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_colour_lookup_table_s1                                 (pipeline_bridge_m1_granted_colour_lookup_table_s1),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_colour_lookup_table_s1                       (pipeline_bridge_m1_qualified_request_colour_lookup_table_s1),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1                         (pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_requests_colour_lookup_table_s1                                (pipeline_bridge_m1_requests_colour_lookup_table_s1),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  colour_lookup_table_s2_arbitrator the_colour_lookup_table_s2
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported                 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_flush_qualified_exported),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_granted_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter                          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_latency_counter),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_qualified_request_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read                                     (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2   (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_read_data_valid_colour_lookup_table_s2),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource0_requests_colour_lookup_table_s2),
      .clk                                                                                                                                                                    (system_clk),
      .colour_lookup_table_s2_address                                                                                                                                         (colour_lookup_table_s2_address),
      .colour_lookup_table_s2_byteenable                                                                                                                                      (colour_lookup_table_s2_byteenable),
      .colour_lookup_table_s2_chipselect                                                                                                                                      (colour_lookup_table_s2_chipselect),
      .colour_lookup_table_s2_clken                                                                                                                                           (colour_lookup_table_s2_clken),
      .colour_lookup_table_s2_readdata                                                                                                                                        (colour_lookup_table_s2_readdata),
      .colour_lookup_table_s2_readdata_from_sa                                                                                                                                (colour_lookup_table_s2_readdata_from_sa),
      .colour_lookup_table_s2_reset                                                                                                                                           (colour_lookup_table_s2_reset),
      .colour_lookup_table_s2_write                                                                                                                                           (colour_lookup_table_s2_write),
      .colour_lookup_table_s2_writedata                                                                                                                                       (colour_lookup_table_s2_writedata),
      .d1_colour_lookup_table_s2_end_xfer                                                                                                                                     (d1_colour_lookup_table_s2_end_xfer),
      .dummy_master_inst_granted_colour_lookup_table_s2                                                                                                                       (dummy_master_inst_granted_colour_lookup_table_s2),
      .dummy_master_inst_m0_address_to_slave                                                                                                                                  (dummy_master_inst_m0_address_to_slave),
      .dummy_master_inst_m0_write                                                                                                                                             (dummy_master_inst_m0_write),
      .dummy_master_inst_m0_writedata                                                                                                                                         (dummy_master_inst_m0_writedata),
      .dummy_master_inst_qualified_request_colour_lookup_table_s2                                                                                                             (dummy_master_inst_qualified_request_colour_lookup_table_s2),
      .dummy_master_inst_requests_colour_lookup_table_s2                                                                                                                      (dummy_master_inst_requests_colour_lookup_table_s2),
      .reset_n                                                                                                                                                                (system_clk_reset_n)
    );

  colour_lookup_table the_colour_lookup_table
    (
      .address     (colour_lookup_table_s1_address),
      .address2    (colour_lookup_table_s2_address),
      .byteenable  (colour_lookup_table_s1_byteenable),
      .byteenable2 (colour_lookup_table_s2_byteenable),
      .chipselect  (colour_lookup_table_s1_chipselect),
      .chipselect2 (colour_lookup_table_s2_chipselect),
      .clk         (system_clk),
      .clk2        (system_clk),
      .clken       (colour_lookup_table_s1_clken),
      .clken2      (colour_lookup_table_s2_clken),
      .readdata    (colour_lookup_table_s1_readdata),
      .readdata2   (colour_lookup_table_s2_readdata),
      .reset       (colour_lookup_table_s1_reset),
      .reset2      (colour_lookup_table_s2_reset),
      .write       (colour_lookup_table_s1_write),
      .write2      (colour_lookup_table_s2_write),
      .writedata   (colour_lookup_table_s1_writedata),
      .writedata2  (colour_lookup_table_s2_writedata)
    );

  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                                               (system_clk),
      .cpu_jtag_debug_module_address                                                     (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                                               (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                                                  (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                                                  (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                                                 (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                                                    (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                                            (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset_n                                                     (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                                                (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                                        (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                                       (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                                                   (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                                                 (d1_cpu_jtag_debug_module_end_xfer),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                     (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_debugaccess                                                    (pipeline_bridge_m1_debugaccess),
      .pipeline_bridge_m1_granted_cpu_jtag_debug_module                                  (pipeline_bridge_m1_granted_cpu_jtag_debug_module),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module                        (pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module                          (pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_requests_cpu_jtag_debug_module                                 (pipeline_bridge_m1_requests_cpu_jtag_debug_module),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa                       (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_irq_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_readdata_from_sa),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_waitrequest_n_from_sa),
      .clk                                                                                                             (system_clk),
      .cpu_data_master_address                                                                                         (cpu_data_master_address),
      .cpu_data_master_address_to_slave                                                                                (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                                                      (cpu_data_master_byteenable),
      .cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0           (cpu_data_master_granted_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_granted_pipeline_bridge_s1                                                                      (cpu_data_master_granted_pipeline_bridge_s1),
      .cpu_data_master_irq                                                                                             (cpu_data_master_irq),
      .cpu_data_master_latency_counter                                                                                 (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0 (cpu_data_master_qualified_request_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_qualified_request_pipeline_bridge_s1                                                            (cpu_data_master_qualified_request_pipeline_bridge_s1),
      .cpu_data_master_read                                                                                            (cpu_data_master_read),
      .cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0   (cpu_data_master_read_data_valid_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_read_data_valid_pipeline_bridge_s1                                                              (cpu_data_master_read_data_valid_pipeline_bridge_s1),
      .cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register                                               (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register),
      .cpu_data_master_readdata                                                                                        (cpu_data_master_readdata),
      .cpu_data_master_readdatavalid                                                                                   (cpu_data_master_readdatavalid),
      .cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0          (cpu_data_master_requests_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0),
      .cpu_data_master_requests_pipeline_bridge_s1                                                                     (cpu_data_master_requests_pipeline_bridge_s1),
      .cpu_data_master_waitrequest                                                                                     (cpu_data_master_waitrequest),
      .cpu_data_master_write                                                                                           (cpu_data_master_write),
      .cpu_data_master_writedata                                                                                       (cpu_data_master_writedata),
      .d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer                       (d1_accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_cpu_interface0_end_xfer),
      .d1_pipeline_bridge_s1_end_xfer                                                                                  (d1_pipeline_bridge_s1_end_xfer),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                                                         (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .lcd_sgdma_csr_irq_from_sa                                                                                       (lcd_sgdma_csr_irq_from_sa),
      .pipeline_bridge_s1_readdata_from_sa                                                                             (pipeline_bridge_s1_readdata_from_sa),
      .pipeline_bridge_s1_waitrequest_from_sa                                                                          (pipeline_bridge_s1_waitrequest_from_sa),
      .push_buttons_s1_irq_from_sa                                                                                     (push_buttons_s1_irq_from_sa),
      .reset_n                                                                                                         (system_clk_reset_n),
      .system_clk                                                                                                      (system_clk),
      .system_clk_reset_n                                                                                              (system_clk_reset_n),
      .system_tick_s1_irq_from_sa                                                                                      (system_tick_s1_irq_from_sa),
      .touchPanel_irq_n_s1_irq_from_sa                                                                                 (touchPanel_irq_n_s1_irq_from_sa),
      .touchPanel_spi_spi_control_port_irq_from_sa                                                                     (touchPanel_spi_spi_control_port_irq_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                                      (system_clk),
      .cpu_instruction_master_address                                           (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                                  (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_pipeline_bridge_s1                        (cpu_instruction_master_granted_pipeline_bridge_s1),
      .cpu_instruction_master_latency_counter                                   (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_pipeline_bridge_s1              (cpu_instruction_master_qualified_request_pipeline_bridge_s1),
      .cpu_instruction_master_read                                              (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_s1                (cpu_instruction_master_read_data_valid_pipeline_bridge_s1),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register (cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register),
      .cpu_instruction_master_readdata                                          (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                                     (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_pipeline_bridge_s1                       (cpu_instruction_master_requests_pipeline_bridge_s1),
      .cpu_instruction_master_waitrequest                                       (cpu_instruction_master_waitrequest),
      .d1_pipeline_bridge_s1_end_xfer                                           (d1_pipeline_bridge_s1_end_xfer),
      .pipeline_bridge_s1_readdata_from_sa                                      (pipeline_bridge_s1_readdata_from_sa),
      .pipeline_bridge_s1_waitrequest_from_sa                                   (pipeline_bridge_s1_waitrequest_from_sa),
      .reset_n                                                                  (system_clk_reset_n)
    );

  cpu the_cpu
    (
      .clk                                   (system_clk),
      .d_address                             (cpu_data_master_address),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_readdatavalid                       (cpu_data_master_readdatavalid),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  ddr_sdram_clock_crossing_bridge_s1_arbitrator the_ddr_sdram_clock_crossing_bridge_s1
    (
      .clk                                                                                               (system_clk),
      .d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer                                                    (d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer),
      .ddr_sdram_clock_crossing_bridge_s1_address                                                        (ddr_sdram_clock_crossing_bridge_s1_address),
      .ddr_sdram_clock_crossing_bridge_s1_byteenable                                                     (ddr_sdram_clock_crossing_bridge_s1_byteenable),
      .ddr_sdram_clock_crossing_bridge_s1_endofpacket                                                    (ddr_sdram_clock_crossing_bridge_s1_endofpacket),
      .ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa                                            (ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa),
      .ddr_sdram_clock_crossing_bridge_s1_nativeaddress                                                  (ddr_sdram_clock_crossing_bridge_s1_nativeaddress),
      .ddr_sdram_clock_crossing_bridge_s1_read                                                           (ddr_sdram_clock_crossing_bridge_s1_read),
      .ddr_sdram_clock_crossing_bridge_s1_readdata                                                       (ddr_sdram_clock_crossing_bridge_s1_readdata),
      .ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa                                               (ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa),
      .ddr_sdram_clock_crossing_bridge_s1_readdatavalid                                                  (ddr_sdram_clock_crossing_bridge_s1_readdatavalid),
      .ddr_sdram_clock_crossing_bridge_s1_reset_n                                                        (ddr_sdram_clock_crossing_bridge_s1_reset_n),
      .ddr_sdram_clock_crossing_bridge_s1_waitrequest                                                    (ddr_sdram_clock_crossing_bridge_s1_waitrequest),
      .ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa                                            (ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa),
      .ddr_sdram_clock_crossing_bridge_s1_write                                                          (ddr_sdram_clock_crossing_bridge_s1_write),
      .ddr_sdram_clock_crossing_bridge_s1_writedata                                                      (ddr_sdram_clock_crossing_bridge_s1_writedata),
      .frame_buffer_pipeline_bridge_m1_address_to_slave                                                  (frame_buffer_pipeline_bridge_m1_address_to_slave),
      .frame_buffer_pipeline_bridge_m1_burstcount                                                        (frame_buffer_pipeline_bridge_m1_burstcount),
      .frame_buffer_pipeline_bridge_m1_byteenable                                                        (frame_buffer_pipeline_bridge_m1_byteenable),
      .frame_buffer_pipeline_bridge_m1_chipselect                                                        (frame_buffer_pipeline_bridge_m1_chipselect),
      .frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1                        (frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_latency_counter                                                   (frame_buffer_pipeline_bridge_m1_latency_counter),
      .frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1              (frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_read                                                              (frame_buffer_pipeline_bridge_m1_read),
      .frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1                (frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register (frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register),
      .frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1                       (frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_write                                                             (frame_buffer_pipeline_bridge_m1_write),
      .frame_buffer_pipeline_bridge_m1_writedata                                                         (frame_buffer_pipeline_bridge_m1_writedata),
      .reset_n                                                                                           (system_clk_reset_n)
    );

  ddr_sdram_clock_crossing_bridge_m1_arbitrator the_ddr_sdram_clock_crossing_bridge_m1
    (
      .clk                                                                               (frame_buffer_phy_clk_out),
      .d1_frame_buffer_s1_end_xfer                                                       (d1_frame_buffer_s1_end_xfer),
      .ddr_sdram_clock_crossing_bridge_m1_address                                        (ddr_sdram_clock_crossing_bridge_m1_address),
      .ddr_sdram_clock_crossing_bridge_m1_address_to_slave                               (ddr_sdram_clock_crossing_bridge_m1_address_to_slave),
      .ddr_sdram_clock_crossing_bridge_m1_byteenable                                     (ddr_sdram_clock_crossing_bridge_m1_byteenable),
      .ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1                        (ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_latency_counter                                (ddr_sdram_clock_crossing_bridge_m1_latency_counter),
      .ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1              (ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_read                                           (ddr_sdram_clock_crossing_bridge_m1_read),
      .ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1                (ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register (ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register),
      .ddr_sdram_clock_crossing_bridge_m1_readdata                                       (ddr_sdram_clock_crossing_bridge_m1_readdata),
      .ddr_sdram_clock_crossing_bridge_m1_readdatavalid                                  (ddr_sdram_clock_crossing_bridge_m1_readdatavalid),
      .ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1                       (ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_reset_n                                        (ddr_sdram_clock_crossing_bridge_m1_reset_n),
      .ddr_sdram_clock_crossing_bridge_m1_waitrequest                                    (ddr_sdram_clock_crossing_bridge_m1_waitrequest),
      .ddr_sdram_clock_crossing_bridge_m1_write                                          (ddr_sdram_clock_crossing_bridge_m1_write),
      .ddr_sdram_clock_crossing_bridge_m1_writedata                                      (ddr_sdram_clock_crossing_bridge_m1_writedata),
      .frame_buffer_s1_readdata_from_sa                                                  (frame_buffer_s1_readdata_from_sa),
      .frame_buffer_s1_waitrequest_n_from_sa                                             (frame_buffer_s1_waitrequest_n_from_sa),
      .reset_n                                                                           (frame_buffer_phy_clk_out_reset_n)
    );

  ddr_sdram_clock_crossing_bridge the_ddr_sdram_clock_crossing_bridge
    (
      .master_address       (ddr_sdram_clock_crossing_bridge_m1_address),
      .master_byteenable    (ddr_sdram_clock_crossing_bridge_m1_byteenable),
      .master_clk           (frame_buffer_phy_clk_out),
      .master_endofpacket   (ddr_sdram_clock_crossing_bridge_m1_endofpacket),
      .master_nativeaddress (ddr_sdram_clock_crossing_bridge_m1_nativeaddress),
      .master_read          (ddr_sdram_clock_crossing_bridge_m1_read),
      .master_readdata      (ddr_sdram_clock_crossing_bridge_m1_readdata),
      .master_readdatavalid (ddr_sdram_clock_crossing_bridge_m1_readdatavalid),
      .master_reset_n       (ddr_sdram_clock_crossing_bridge_m1_reset_n),
      .master_waitrequest   (ddr_sdram_clock_crossing_bridge_m1_waitrequest),
      .master_write         (ddr_sdram_clock_crossing_bridge_m1_write),
      .master_writedata     (ddr_sdram_clock_crossing_bridge_m1_writedata),
      .slave_address        (ddr_sdram_clock_crossing_bridge_s1_address),
      .slave_byteenable     (ddr_sdram_clock_crossing_bridge_s1_byteenable),
      .slave_clk            (system_clk),
      .slave_endofpacket    (ddr_sdram_clock_crossing_bridge_s1_endofpacket),
      .slave_nativeaddress  (ddr_sdram_clock_crossing_bridge_s1_nativeaddress),
      .slave_read           (ddr_sdram_clock_crossing_bridge_s1_read),
      .slave_readdata       (ddr_sdram_clock_crossing_bridge_s1_readdata),
      .slave_readdatavalid  (ddr_sdram_clock_crossing_bridge_s1_readdatavalid),
      .slave_reset_n        (ddr_sdram_clock_crossing_bridge_s1_reset_n),
      .slave_waitrequest    (ddr_sdram_clock_crossing_bridge_s1_waitrequest),
      .slave_write          (ddr_sdram_clock_crossing_bridge_s1_write),
      .slave_writedata      (ddr_sdram_clock_crossing_bridge_s1_writedata)
    );

  descriptor_memory_s1_arbitrator the_descriptor_memory_s1
    (
      .clk                                                                               (system_clk),
      .d1_descriptor_memory_s1_end_xfer                                                  (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_address                                                      (descriptor_memory_s1_address),
      .descriptor_memory_s1_byteenable                                                   (descriptor_memory_s1_byteenable),
      .descriptor_memory_s1_chipselect                                                   (descriptor_memory_s1_chipselect),
      .descriptor_memory_s1_clken                                                        (descriptor_memory_s1_clken),
      .descriptor_memory_s1_readdata                                                     (descriptor_memory_s1_readdata),
      .descriptor_memory_s1_readdata_from_sa                                             (descriptor_memory_s1_readdata_from_sa),
      .descriptor_memory_s1_reset                                                        (descriptor_memory_s1_reset),
      .descriptor_memory_s1_write                                                        (descriptor_memory_s1_write),
      .descriptor_memory_s1_writedata                                                    (descriptor_memory_s1_writedata),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                     (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_descriptor_memory_s1                                   (pipeline_bridge_m1_granted_descriptor_memory_s1),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_descriptor_memory_s1                         (pipeline_bridge_m1_qualified_request_descriptor_memory_s1),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_descriptor_memory_s1                           (pipeline_bridge_m1_read_data_valid_descriptor_memory_s1),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_requests_descriptor_memory_s1                                  (pipeline_bridge_m1_requests_descriptor_memory_s1),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  descriptor_memory_s2_arbitrator the_descriptor_memory_s2
    (
      .clk                                                               (system_clk),
      .d1_descriptor_memory_s2_end_xfer                                  (d1_descriptor_memory_s2_end_xfer),
      .descriptor_memory_s2_address                                      (descriptor_memory_s2_address),
      .descriptor_memory_s2_byteenable                                   (descriptor_memory_s2_byteenable),
      .descriptor_memory_s2_chipselect                                   (descriptor_memory_s2_chipselect),
      .descriptor_memory_s2_clken                                        (descriptor_memory_s2_clken),
      .descriptor_memory_s2_readdata                                     (descriptor_memory_s2_readdata),
      .descriptor_memory_s2_readdata_from_sa                             (descriptor_memory_s2_readdata_from_sa),
      .descriptor_memory_s2_reset                                        (descriptor_memory_s2_reset),
      .descriptor_memory_s2_write                                        (descriptor_memory_s2_write),
      .descriptor_memory_s2_writedata                                    (descriptor_memory_s2_writedata),
      .lcd_sgdma_descriptor_read_address_to_slave                        (lcd_sgdma_descriptor_read_address_to_slave),
      .lcd_sgdma_descriptor_read_granted_descriptor_memory_s2            (lcd_sgdma_descriptor_read_granted_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_latency_counter                         (lcd_sgdma_descriptor_read_latency_counter),
      .lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2  (lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_read                                    (lcd_sgdma_descriptor_read_read),
      .lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2    (lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_requests_descriptor_memory_s2           (lcd_sgdma_descriptor_read_requests_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_address_to_slave                       (lcd_sgdma_descriptor_write_address_to_slave),
      .lcd_sgdma_descriptor_write_granted_descriptor_memory_s2           (lcd_sgdma_descriptor_write_granted_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2 (lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_requests_descriptor_memory_s2          (lcd_sgdma_descriptor_write_requests_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_write                                  (lcd_sgdma_descriptor_write_write),
      .lcd_sgdma_descriptor_write_writedata                              (lcd_sgdma_descriptor_write_writedata),
      .reset_n                                                           (system_clk_reset_n)
    );

  descriptor_memory the_descriptor_memory
    (
      .address     (descriptor_memory_s1_address),
      .address2    (descriptor_memory_s2_address),
      .byteenable  (descriptor_memory_s1_byteenable),
      .byteenable2 (descriptor_memory_s2_byteenable),
      .chipselect  (descriptor_memory_s1_chipselect),
      .chipselect2 (descriptor_memory_s2_chipselect),
      .clk         (system_clk),
      .clk2        (system_clk),
      .clken       (descriptor_memory_s1_clken),
      .clken2      (descriptor_memory_s2_clken),
      .readdata    (descriptor_memory_s1_readdata),
      .readdata2   (descriptor_memory_s2_readdata),
      .reset       (descriptor_memory_s1_reset),
      .reset2      (descriptor_memory_s2_reset),
      .write       (descriptor_memory_s1_write),
      .write2      (descriptor_memory_s2_write),
      .writedata   (descriptor_memory_s1_writedata),
      .writedata2  (descriptor_memory_s2_writedata)
    );

  dummy_master_inst_m0_arbitrator the_dummy_master_inst_m0
    (
      .clk                                                        (system_clk),
      .d1_colour_lookup_table_s2_end_xfer                         (d1_colour_lookup_table_s2_end_xfer),
      .dummy_master_inst_granted_colour_lookup_table_s2           (dummy_master_inst_granted_colour_lookup_table_s2),
      .dummy_master_inst_m0_address                               (dummy_master_inst_m0_address),
      .dummy_master_inst_m0_address_to_slave                      (dummy_master_inst_m0_address_to_slave),
      .dummy_master_inst_m0_waitrequest                           (dummy_master_inst_m0_waitrequest),
      .dummy_master_inst_m0_write                                 (dummy_master_inst_m0_write),
      .dummy_master_inst_m0_writedata                             (dummy_master_inst_m0_writedata),
      .dummy_master_inst_qualified_request_colour_lookup_table_s2 (dummy_master_inst_qualified_request_colour_lookup_table_s2),
      .dummy_master_inst_requests_colour_lookup_table_s2          (dummy_master_inst_requests_colour_lookup_table_s2),
      .reset_n                                                    (system_clk_reset_n)
    );

  dummy_master_inst the_dummy_master_inst
    (
      .address     (dummy_master_inst_m0_address),
      .waitrequest (dummy_master_inst_m0_waitrequest),
      .write       (dummy_master_inst_m0_write),
      .writedata   (dummy_master_inst_m0_writedata)
    );

  flash_ssram_pipeline_bridge_s1_arbitrator the_flash_ssram_pipeline_bridge_s1
    (
      .clk                                                                               (system_clk),
      .d1_flash_ssram_pipeline_bridge_s1_end_xfer                                        (d1_flash_ssram_pipeline_bridge_s1_end_xfer),
      .flash_ssram_pipeline_bridge_s1_address                                            (flash_ssram_pipeline_bridge_s1_address),
      .flash_ssram_pipeline_bridge_s1_arbiterlock                                        (flash_ssram_pipeline_bridge_s1_arbiterlock),
      .flash_ssram_pipeline_bridge_s1_arbiterlock2                                       (flash_ssram_pipeline_bridge_s1_arbiterlock2),
      .flash_ssram_pipeline_bridge_s1_burstcount                                         (flash_ssram_pipeline_bridge_s1_burstcount),
      .flash_ssram_pipeline_bridge_s1_byteenable                                         (flash_ssram_pipeline_bridge_s1_byteenable),
      .flash_ssram_pipeline_bridge_s1_chipselect                                         (flash_ssram_pipeline_bridge_s1_chipselect),
      .flash_ssram_pipeline_bridge_s1_debugaccess                                        (flash_ssram_pipeline_bridge_s1_debugaccess),
      .flash_ssram_pipeline_bridge_s1_endofpacket                                        (flash_ssram_pipeline_bridge_s1_endofpacket),
      .flash_ssram_pipeline_bridge_s1_endofpacket_from_sa                                (flash_ssram_pipeline_bridge_s1_endofpacket_from_sa),
      .flash_ssram_pipeline_bridge_s1_nativeaddress                                      (flash_ssram_pipeline_bridge_s1_nativeaddress),
      .flash_ssram_pipeline_bridge_s1_read                                               (flash_ssram_pipeline_bridge_s1_read),
      .flash_ssram_pipeline_bridge_s1_readdata                                           (flash_ssram_pipeline_bridge_s1_readdata),
      .flash_ssram_pipeline_bridge_s1_readdata_from_sa                                   (flash_ssram_pipeline_bridge_s1_readdata_from_sa),
      .flash_ssram_pipeline_bridge_s1_readdatavalid                                      (flash_ssram_pipeline_bridge_s1_readdatavalid),
      .flash_ssram_pipeline_bridge_s1_reset_n                                            (flash_ssram_pipeline_bridge_s1_reset_n),
      .flash_ssram_pipeline_bridge_s1_waitrequest                                        (flash_ssram_pipeline_bridge_s1_waitrequest),
      .flash_ssram_pipeline_bridge_s1_waitrequest_from_sa                                (flash_ssram_pipeline_bridge_s1_waitrequest_from_sa),
      .flash_ssram_pipeline_bridge_s1_write                                              (flash_ssram_pipeline_bridge_s1_write),
      .flash_ssram_pipeline_bridge_s1_writedata                                          (flash_ssram_pipeline_bridge_s1_writedata),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                     (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_debugaccess                                                    (pipeline_bridge_m1_debugaccess),
      .pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1                         (pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1               (pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1                 (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1                        (pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  flash_ssram_pipeline_bridge_m1_arbitrator the_flash_ssram_pipeline_bridge_m1
    (
      .clk                                                       (system_clk),
      .d1_tristate_bridge_avalon_slave_end_xfer                  (d1_tristate_bridge_avalon_slave_end_xfer),
      .flash_s1_wait_counter_eq_0                                (flash_s1_wait_counter_eq_0),
      .flash_ssram_pipeline_bridge_m1_address                    (flash_ssram_pipeline_bridge_m1_address),
      .flash_ssram_pipeline_bridge_m1_address_to_slave           (flash_ssram_pipeline_bridge_m1_address_to_slave),
      .flash_ssram_pipeline_bridge_m1_burstcount                 (flash_ssram_pipeline_bridge_m1_burstcount),
      .flash_ssram_pipeline_bridge_m1_byteenable                 (flash_ssram_pipeline_bridge_m1_byteenable),
      .flash_ssram_pipeline_bridge_m1_byteenable_flash_s1        (flash_ssram_pipeline_bridge_m1_byteenable_flash_s1),
      .flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1        (flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_chipselect                 (flash_ssram_pipeline_bridge_m1_chipselect),
      .flash_ssram_pipeline_bridge_m1_dbs_address                (flash_ssram_pipeline_bridge_m1_dbs_address),
      .flash_ssram_pipeline_bridge_m1_dbs_write_16               (flash_ssram_pipeline_bridge_m1_dbs_write_16),
      .flash_ssram_pipeline_bridge_m1_dbs_write_32               (flash_ssram_pipeline_bridge_m1_dbs_write_32),
      .flash_ssram_pipeline_bridge_m1_granted_flash_s1           (flash_ssram_pipeline_bridge_m1_granted_flash_s1),
      .flash_ssram_pipeline_bridge_m1_granted_ssram_s1           (flash_ssram_pipeline_bridge_m1_granted_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_latency_counter            (flash_ssram_pipeline_bridge_m1_latency_counter),
      .flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 (flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1),
      .flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1 (flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_read                       (flash_ssram_pipeline_bridge_m1_read),
      .flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1   (flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1),
      .flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1   (flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_readdata                   (flash_ssram_pipeline_bridge_m1_readdata),
      .flash_ssram_pipeline_bridge_m1_readdatavalid              (flash_ssram_pipeline_bridge_m1_readdatavalid),
      .flash_ssram_pipeline_bridge_m1_requests_flash_s1          (flash_ssram_pipeline_bridge_m1_requests_flash_s1),
      .flash_ssram_pipeline_bridge_m1_requests_ssram_s1          (flash_ssram_pipeline_bridge_m1_requests_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_waitrequest                (flash_ssram_pipeline_bridge_m1_waitrequest),
      .flash_ssram_pipeline_bridge_m1_write                      (flash_ssram_pipeline_bridge_m1_write),
      .flash_ssram_pipeline_bridge_m1_writedata                  (flash_ssram_pipeline_bridge_m1_writedata),
      .incoming_tristate_bridge_data                             (incoming_tristate_bridge_data),
      .incoming_tristate_bridge_data_with_Xs_converted_to_0      (incoming_tristate_bridge_data_with_Xs_converted_to_0),
      .reset_n                                                   (system_clk_reset_n)
    );

  flash_ssram_pipeline_bridge the_flash_ssram_pipeline_bridge
    (
      .clk              (system_clk),
      .m1_address       (flash_ssram_pipeline_bridge_m1_address),
      .m1_burstcount    (flash_ssram_pipeline_bridge_m1_burstcount),
      .m1_byteenable    (flash_ssram_pipeline_bridge_m1_byteenable),
      .m1_chipselect    (flash_ssram_pipeline_bridge_m1_chipselect),
      .m1_debugaccess   (flash_ssram_pipeline_bridge_m1_debugaccess),
      .m1_endofpacket   (flash_ssram_pipeline_bridge_m1_endofpacket),
      .m1_read          (flash_ssram_pipeline_bridge_m1_read),
      .m1_readdata      (flash_ssram_pipeline_bridge_m1_readdata),
      .m1_readdatavalid (flash_ssram_pipeline_bridge_m1_readdatavalid),
      .m1_waitrequest   (flash_ssram_pipeline_bridge_m1_waitrequest),
      .m1_write         (flash_ssram_pipeline_bridge_m1_write),
      .m1_writedata     (flash_ssram_pipeline_bridge_m1_writedata),
      .reset_n          (flash_ssram_pipeline_bridge_s1_reset_n),
      .s1_address       (flash_ssram_pipeline_bridge_s1_address),
      .s1_arbiterlock   (flash_ssram_pipeline_bridge_s1_arbiterlock),
      .s1_arbiterlock2  (flash_ssram_pipeline_bridge_s1_arbiterlock2),
      .s1_burstcount    (flash_ssram_pipeline_bridge_s1_burstcount),
      .s1_byteenable    (flash_ssram_pipeline_bridge_s1_byteenable),
      .s1_chipselect    (flash_ssram_pipeline_bridge_s1_chipselect),
      .s1_debugaccess   (flash_ssram_pipeline_bridge_s1_debugaccess),
      .s1_endofpacket   (flash_ssram_pipeline_bridge_s1_endofpacket),
      .s1_nativeaddress (flash_ssram_pipeline_bridge_s1_nativeaddress),
      .s1_read          (flash_ssram_pipeline_bridge_s1_read),
      .s1_readdata      (flash_ssram_pipeline_bridge_s1_readdata),
      .s1_readdatavalid (flash_ssram_pipeline_bridge_s1_readdatavalid),
      .s1_waitrequest   (flash_ssram_pipeline_bridge_s1_waitrequest),
      .s1_write         (flash_ssram_pipeline_bridge_s1_write),
      .s1_writedata     (flash_ssram_pipeline_bridge_s1_writedata)
    );

  frame_buffer_s1_arbitrator the_frame_buffer_s1
    (
      .clk                                                                               (frame_buffer_phy_clk_out),
      .d1_frame_buffer_s1_end_xfer                                                       (d1_frame_buffer_s1_end_xfer),
      .ddr_sdram_clock_crossing_bridge_m1_address_to_slave                               (ddr_sdram_clock_crossing_bridge_m1_address_to_slave),
      .ddr_sdram_clock_crossing_bridge_m1_byteenable                                     (ddr_sdram_clock_crossing_bridge_m1_byteenable),
      .ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1                        (ddr_sdram_clock_crossing_bridge_m1_granted_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_latency_counter                                (ddr_sdram_clock_crossing_bridge_m1_latency_counter),
      .ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1              (ddr_sdram_clock_crossing_bridge_m1_qualified_request_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_read                                           (ddr_sdram_clock_crossing_bridge_m1_read),
      .ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1                (ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register (ddr_sdram_clock_crossing_bridge_m1_read_data_valid_frame_buffer_s1_shift_register),
      .ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1                       (ddr_sdram_clock_crossing_bridge_m1_requests_frame_buffer_s1),
      .ddr_sdram_clock_crossing_bridge_m1_write                                          (ddr_sdram_clock_crossing_bridge_m1_write),
      .ddr_sdram_clock_crossing_bridge_m1_writedata                                      (ddr_sdram_clock_crossing_bridge_m1_writedata),
      .frame_buffer_s1_address                                                           (frame_buffer_s1_address),
      .frame_buffer_s1_beginbursttransfer                                                (frame_buffer_s1_beginbursttransfer),
      .frame_buffer_s1_burstcount                                                        (frame_buffer_s1_burstcount),
      .frame_buffer_s1_byteenable                                                        (frame_buffer_s1_byteenable),
      .frame_buffer_s1_read                                                              (frame_buffer_s1_read),
      .frame_buffer_s1_readdata                                                          (frame_buffer_s1_readdata),
      .frame_buffer_s1_readdata_from_sa                                                  (frame_buffer_s1_readdata_from_sa),
      .frame_buffer_s1_readdatavalid                                                     (frame_buffer_s1_readdatavalid),
      .frame_buffer_s1_resetrequest_n                                                    (frame_buffer_s1_resetrequest_n),
      .frame_buffer_s1_resetrequest_n_from_sa                                            (frame_buffer_s1_resetrequest_n_from_sa),
      .frame_buffer_s1_waitrequest_n                                                     (frame_buffer_s1_waitrequest_n),
      .frame_buffer_s1_waitrequest_n_from_sa                                             (frame_buffer_s1_waitrequest_n_from_sa),
      .frame_buffer_s1_write                                                             (frame_buffer_s1_write),
      .frame_buffer_s1_writedata                                                         (frame_buffer_s1_writedata),
      .reset_n                                                                           (frame_buffer_phy_clk_out_reset_n)
    );

  //frame_buffer_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  assign frame_buffer_aux_full_rate_clk_out = out_clk_frame_buffer_aux_full_rate_clk;

  //frame_buffer_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  assign frame_buffer_aux_half_rate_clk_out = out_clk_frame_buffer_aux_half_rate_clk;

  //frame_buffer_phy_clk_out out_clk assignment, which is an e_assign
  assign frame_buffer_phy_clk_out = out_clk_frame_buffer_phy_clk;

  //reset is asserted asynchronously and deasserted synchronously
  system_reset_ext_clk_one_domain_synch_module system_reset_ext_clk_one_domain_synch
    (
      .clk      (ext_clk_one),
      .data_in  (1'b1),
      .data_out (ext_clk_one_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa |
    0 |
    ~frame_buffer_s1_resetrequest_n_from_sa |
    ~frame_buffer_s1_resetrequest_n_from_sa |
    0 |
    0);

  frame_buffer the_frame_buffer
    (
      .aux_full_rate_clk (out_clk_frame_buffer_aux_full_rate_clk),
      .aux_half_rate_clk (out_clk_frame_buffer_aux_half_rate_clk),
      .global_reset_n    (global_reset_n_to_the_frame_buffer),
      .local_address     (frame_buffer_s1_address),
      .local_be          (frame_buffer_s1_byteenable),
      .local_burstbegin  (frame_buffer_s1_beginbursttransfer),
      .local_init_done   (local_init_done_from_the_frame_buffer),
      .local_rdata       (frame_buffer_s1_readdata),
      .local_rdata_valid (frame_buffer_s1_readdatavalid),
      .local_read_req    (frame_buffer_s1_read),
      .local_ready       (frame_buffer_s1_waitrequest_n),
      .local_refresh_ack (local_refresh_ack_from_the_frame_buffer),
      .local_size        (frame_buffer_s1_burstcount),
      .local_wdata       (frame_buffer_s1_writedata),
      .local_wdata_req   (local_wdata_req_from_the_frame_buffer),
      .local_write_req   (frame_buffer_s1_write),
      .mem_addr          (mem_addr_from_the_frame_buffer),
      .mem_ba            (mem_ba_from_the_frame_buffer),
      .mem_cas_n         (mem_cas_n_from_the_frame_buffer),
      .mem_cke           (mem_cke_from_the_frame_buffer),
      .mem_clk           (mem_clk_to_and_from_the_frame_buffer),
      .mem_clk_n         (mem_clk_n_to_and_from_the_frame_buffer),
      .mem_cs_n          (mem_cs_n_from_the_frame_buffer),
      .mem_dm            (mem_dm_from_the_frame_buffer),
      .mem_dq            (mem_dq_to_and_from_the_frame_buffer),
      .mem_dqs           (mem_dqs_to_and_from_the_frame_buffer),
      .mem_ras_n         (mem_ras_n_from_the_frame_buffer),
      .mem_we_n          (mem_we_n_from_the_frame_buffer),
      .phy_clk           (out_clk_frame_buffer_phy_clk),
      .pll_ref_clk       (ext_clk_one),
      .reset_phy_clk_n   (reset_phy_clk_n_from_the_frame_buffer),
      .reset_request_n   (frame_buffer_s1_resetrequest_n),
      .soft_reset_n      (ext_clk_one_reset_n)
    );

  frame_buffer_pipeline_bridge_s1_arbitrator the_frame_buffer_pipeline_bridge_s1
    (
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave                                  (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_address_to_slave),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable                                        (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_byteenable),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1           (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_granted_frame_buffer_pipeline_bridge_s1),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1 (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_qualified_request_frame_buffer_pipeline_bridge_s1),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1          (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_requests_frame_buffer_pipeline_bridge_s1),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write                                             (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_write),
      .accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata                                         (accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_accelerator_mandelbrot_hw_draw_int_mandelbrot_master_resource1_writedata),
      .clk                                                                                                                                                                             (system_clk),
      .d1_frame_buffer_pipeline_bridge_s1_end_xfer                                                                                                                                     (d1_frame_buffer_pipeline_bridge_s1_end_xfer),
      .frame_buffer_pipeline_bridge_s1_address                                                                                                                                         (frame_buffer_pipeline_bridge_s1_address),
      .frame_buffer_pipeline_bridge_s1_arbiterlock                                                                                                                                     (frame_buffer_pipeline_bridge_s1_arbiterlock),
      .frame_buffer_pipeline_bridge_s1_arbiterlock2                                                                                                                                    (frame_buffer_pipeline_bridge_s1_arbiterlock2),
      .frame_buffer_pipeline_bridge_s1_burstcount                                                                                                                                      (frame_buffer_pipeline_bridge_s1_burstcount),
      .frame_buffer_pipeline_bridge_s1_byteenable                                                                                                                                      (frame_buffer_pipeline_bridge_s1_byteenable),
      .frame_buffer_pipeline_bridge_s1_chipselect                                                                                                                                      (frame_buffer_pipeline_bridge_s1_chipselect),
      .frame_buffer_pipeline_bridge_s1_debugaccess                                                                                                                                     (frame_buffer_pipeline_bridge_s1_debugaccess),
      .frame_buffer_pipeline_bridge_s1_endofpacket                                                                                                                                     (frame_buffer_pipeline_bridge_s1_endofpacket),
      .frame_buffer_pipeline_bridge_s1_endofpacket_from_sa                                                                                                                             (frame_buffer_pipeline_bridge_s1_endofpacket_from_sa),
      .frame_buffer_pipeline_bridge_s1_nativeaddress                                                                                                                                   (frame_buffer_pipeline_bridge_s1_nativeaddress),
      .frame_buffer_pipeline_bridge_s1_read                                                                                                                                            (frame_buffer_pipeline_bridge_s1_read),
      .frame_buffer_pipeline_bridge_s1_readdata                                                                                                                                        (frame_buffer_pipeline_bridge_s1_readdata),
      .frame_buffer_pipeline_bridge_s1_readdata_from_sa                                                                                                                                (frame_buffer_pipeline_bridge_s1_readdata_from_sa),
      .frame_buffer_pipeline_bridge_s1_readdatavalid                                                                                                                                   (frame_buffer_pipeline_bridge_s1_readdatavalid),
      .frame_buffer_pipeline_bridge_s1_reset_n                                                                                                                                         (frame_buffer_pipeline_bridge_s1_reset_n),
      .frame_buffer_pipeline_bridge_s1_waitrequest                                                                                                                                     (frame_buffer_pipeline_bridge_s1_waitrequest),
      .frame_buffer_pipeline_bridge_s1_waitrequest_from_sa                                                                                                                             (frame_buffer_pipeline_bridge_s1_waitrequest_from_sa),
      .frame_buffer_pipeline_bridge_s1_write                                                                                                                                           (frame_buffer_pipeline_bridge_s1_write),
      .frame_buffer_pipeline_bridge_s1_writedata                                                                                                                                       (frame_buffer_pipeline_bridge_s1_writedata),
      .lcd_sgdma_m_read_address_to_slave                                                                                                                                               (lcd_sgdma_m_read_address_to_slave),
      .lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1                                                                                                                        (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_latency_counter                                                                                                                                                (lcd_sgdma_m_read_latency_counter),
      .lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1                                                                                                              (lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_read                                                                                                                                                           (lcd_sgdma_m_read_read),
      .lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1                                                                                                                (lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register                                                                                                 (lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1                                                                                                                       (lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_address_to_slave                                                                                                                                             (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                                                                                                                   (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                                                                                                                   (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                                                                                                                   (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_debugaccess                                                                                                                                                  (pipeline_bridge_m1_debugaccess),
      .pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1                                                                                                                      (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_latency_counter                                                                                                                                              (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1                                                                                                            (pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_read                                                                                                                                                         (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register                                                                                                      (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register                                                                                                (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1                                                                                                              (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register                                                                                               (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1                                                                                                                     (pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_write                                                                                                                                                        (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                                                                                                                    (pipeline_bridge_m1_writedata),
      .reset_n                                                                                                                                                                         (system_clk_reset_n)
    );

  frame_buffer_pipeline_bridge_m1_arbitrator the_frame_buffer_pipeline_bridge_m1
    (
      .clk                                                                                               (system_clk),
      .d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer                                                    (d1_ddr_sdram_clock_crossing_bridge_s1_end_xfer),
      .ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa                                            (ddr_sdram_clock_crossing_bridge_s1_endofpacket_from_sa),
      .ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa                                               (ddr_sdram_clock_crossing_bridge_s1_readdata_from_sa),
      .ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa                                            (ddr_sdram_clock_crossing_bridge_s1_waitrequest_from_sa),
      .frame_buffer_pipeline_bridge_m1_address                                                           (frame_buffer_pipeline_bridge_m1_address),
      .frame_buffer_pipeline_bridge_m1_address_to_slave                                                  (frame_buffer_pipeline_bridge_m1_address_to_slave),
      .frame_buffer_pipeline_bridge_m1_burstcount                                                        (frame_buffer_pipeline_bridge_m1_burstcount),
      .frame_buffer_pipeline_bridge_m1_byteenable                                                        (frame_buffer_pipeline_bridge_m1_byteenable),
      .frame_buffer_pipeline_bridge_m1_chipselect                                                        (frame_buffer_pipeline_bridge_m1_chipselect),
      .frame_buffer_pipeline_bridge_m1_endofpacket                                                       (frame_buffer_pipeline_bridge_m1_endofpacket),
      .frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1                        (frame_buffer_pipeline_bridge_m1_granted_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_latency_counter                                                   (frame_buffer_pipeline_bridge_m1_latency_counter),
      .frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1              (frame_buffer_pipeline_bridge_m1_qualified_request_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_read                                                              (frame_buffer_pipeline_bridge_m1_read),
      .frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1                (frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register (frame_buffer_pipeline_bridge_m1_read_data_valid_ddr_sdram_clock_crossing_bridge_s1_shift_register),
      .frame_buffer_pipeline_bridge_m1_readdata                                                          (frame_buffer_pipeline_bridge_m1_readdata),
      .frame_buffer_pipeline_bridge_m1_readdatavalid                                                     (frame_buffer_pipeline_bridge_m1_readdatavalid),
      .frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1                       (frame_buffer_pipeline_bridge_m1_requests_ddr_sdram_clock_crossing_bridge_s1),
      .frame_buffer_pipeline_bridge_m1_waitrequest                                                       (frame_buffer_pipeline_bridge_m1_waitrequest),
      .frame_buffer_pipeline_bridge_m1_write                                                             (frame_buffer_pipeline_bridge_m1_write),
      .frame_buffer_pipeline_bridge_m1_writedata                                                         (frame_buffer_pipeline_bridge_m1_writedata),
      .reset_n                                                                                           (system_clk_reset_n)
    );

  frame_buffer_pipeline_bridge the_frame_buffer_pipeline_bridge
    (
      .clk              (system_clk),
      .m1_address       (frame_buffer_pipeline_bridge_m1_address),
      .m1_burstcount    (frame_buffer_pipeline_bridge_m1_burstcount),
      .m1_byteenable    (frame_buffer_pipeline_bridge_m1_byteenable),
      .m1_chipselect    (frame_buffer_pipeline_bridge_m1_chipselect),
      .m1_debugaccess   (frame_buffer_pipeline_bridge_m1_debugaccess),
      .m1_endofpacket   (frame_buffer_pipeline_bridge_m1_endofpacket),
      .m1_read          (frame_buffer_pipeline_bridge_m1_read),
      .m1_readdata      (frame_buffer_pipeline_bridge_m1_readdata),
      .m1_readdatavalid (frame_buffer_pipeline_bridge_m1_readdatavalid),
      .m1_waitrequest   (frame_buffer_pipeline_bridge_m1_waitrequest),
      .m1_write         (frame_buffer_pipeline_bridge_m1_write),
      .m1_writedata     (frame_buffer_pipeline_bridge_m1_writedata),
      .reset_n          (frame_buffer_pipeline_bridge_s1_reset_n),
      .s1_address       (frame_buffer_pipeline_bridge_s1_address),
      .s1_arbiterlock   (frame_buffer_pipeline_bridge_s1_arbiterlock),
      .s1_arbiterlock2  (frame_buffer_pipeline_bridge_s1_arbiterlock2),
      .s1_burstcount    (frame_buffer_pipeline_bridge_s1_burstcount),
      .s1_byteenable    (frame_buffer_pipeline_bridge_s1_byteenable),
      .s1_chipselect    (frame_buffer_pipeline_bridge_s1_chipselect),
      .s1_debugaccess   (frame_buffer_pipeline_bridge_s1_debugaccess),
      .s1_endofpacket   (frame_buffer_pipeline_bridge_s1_endofpacket),
      .s1_nativeaddress (frame_buffer_pipeline_bridge_s1_nativeaddress),
      .s1_read          (frame_buffer_pipeline_bridge_s1_read),
      .s1_readdata      (frame_buffer_pipeline_bridge_s1_readdata),
      .s1_readdatavalid (frame_buffer_pipeline_bridge_s1_readdatavalid),
      .s1_waitrequest   (frame_buffer_pipeline_bridge_s1_waitrequest),
      .s1_write         (frame_buffer_pipeline_bridge_s1_write),
      .s1_writedata     (frame_buffer_pipeline_bridge_s1_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                                    (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                              (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave           (clock_crossing_bridge_m1_granted_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_latency_counter                               (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                                 (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave (clock_crossing_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_read                                          (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave   (clock_crossing_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave          (clock_crossing_bridge_m1_requests_jtag_uart_avalon_jtag_slave),
      .clock_crossing_bridge_m1_write                                         (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                                     (clock_crossing_bridge_m1_writedata),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                                    (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                                 (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                              (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa                      (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                                        (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                                     (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                                   (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                           (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                               (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa                       (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                                    (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                                (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                        (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                                    (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                                  (jtag_uart_avalon_jtag_slave_writedata),
      .reset_n                                                                (slow_clk_reset_n)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (slow_clk),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  lcd_data_format_adapter_in_arbitrator the_lcd_data_format_adapter_in
    (
      .clk                                      (system_clk),
      .lcd_data_format_adapter_in_data          (lcd_data_format_adapter_in_data),
      .lcd_data_format_adapter_in_empty         (lcd_data_format_adapter_in_empty),
      .lcd_data_format_adapter_in_endofpacket   (lcd_data_format_adapter_in_endofpacket),
      .lcd_data_format_adapter_in_ready         (lcd_data_format_adapter_in_ready),
      .lcd_data_format_adapter_in_ready_from_sa (lcd_data_format_adapter_in_ready_from_sa),
      .lcd_data_format_adapter_in_reset_n       (lcd_data_format_adapter_in_reset_n),
      .lcd_data_format_adapter_in_startofpacket (lcd_data_format_adapter_in_startofpacket),
      .lcd_data_format_adapter_in_valid         (lcd_data_format_adapter_in_valid),
      .lcd_pixel_converter_out_data             (lcd_pixel_converter_out_data),
      .lcd_pixel_converter_out_empty            (lcd_pixel_converter_out_empty),
      .lcd_pixel_converter_out_endofpacket      (lcd_pixel_converter_out_endofpacket),
      .lcd_pixel_converter_out_startofpacket    (lcd_pixel_converter_out_startofpacket),
      .lcd_pixel_converter_out_valid            (lcd_pixel_converter_out_valid),
      .reset_n                                  (system_clk_reset_n)
    );

  lcd_data_format_adapter_out_arbitrator the_lcd_data_format_adapter_out
    (
      .clk                                       (system_clk),
      .lcd_data_format_adapter_out_data          (lcd_data_format_adapter_out_data),
      .lcd_data_format_adapter_out_endofpacket   (lcd_data_format_adapter_out_endofpacket),
      .lcd_data_format_adapter_out_ready         (lcd_data_format_adapter_out_ready),
      .lcd_data_format_adapter_out_startofpacket (lcd_data_format_adapter_out_startofpacket),
      .lcd_data_format_adapter_out_valid         (lcd_data_format_adapter_out_valid),
      .lcd_ta_formatter_to_fifo_in_ready_from_sa (lcd_ta_formatter_to_fifo_in_ready_from_sa),
      .reset_n                                   (system_clk_reset_n)
    );

  lcd_data_format_adapter the_lcd_data_format_adapter
    (
      .clk               (system_clk),
      .in_data           (lcd_data_format_adapter_in_data),
      .in_empty          (lcd_data_format_adapter_in_empty),
      .in_endofpacket    (lcd_data_format_adapter_in_endofpacket),
      .in_ready          (lcd_data_format_adapter_in_ready),
      .in_startofpacket  (lcd_data_format_adapter_in_startofpacket),
      .in_valid          (lcd_data_format_adapter_in_valid),
      .out_data          (lcd_data_format_adapter_out_data),
      .out_endofpacket   (lcd_data_format_adapter_out_endofpacket),
      .out_ready         (lcd_data_format_adapter_out_ready),
      .out_startofpacket (lcd_data_format_adapter_out_startofpacket),
      .out_valid         (lcd_data_format_adapter_out_valid),
      .reset_n           (lcd_data_format_adapter_in_reset_n)
    );

  lcd_data_format_adapter_1_in_arbitrator the_lcd_data_format_adapter_1_in
    (
      .clk                                        (video_clk),
      .lcd_data_format_adapter_1_in_data          (lcd_data_format_adapter_1_in_data),
      .lcd_data_format_adapter_1_in_endofpacket   (lcd_data_format_adapter_1_in_endofpacket),
      .lcd_data_format_adapter_1_in_ready         (lcd_data_format_adapter_1_in_ready),
      .lcd_data_format_adapter_1_in_ready_from_sa (lcd_data_format_adapter_1_in_ready_from_sa),
      .lcd_data_format_adapter_1_in_reset_n       (lcd_data_format_adapter_1_in_reset_n),
      .lcd_data_format_adapter_1_in_startofpacket (lcd_data_format_adapter_1_in_startofpacket),
      .lcd_data_format_adapter_1_in_valid         (lcd_data_format_adapter_1_in_valid),
      .lcd_ta_fifo_to_sequencer_out_data          (lcd_ta_fifo_to_sequencer_out_data),
      .lcd_ta_fifo_to_sequencer_out_endofpacket   (lcd_ta_fifo_to_sequencer_out_endofpacket),
      .lcd_ta_fifo_to_sequencer_out_startofpacket (lcd_ta_fifo_to_sequencer_out_startofpacket),
      .lcd_ta_fifo_to_sequencer_out_valid         (lcd_ta_fifo_to_sequencer_out_valid),
      .reset_n                                    (video_clk_reset_n)
    );

  lcd_data_format_adapter_1_out_arbitrator the_lcd_data_format_adapter_1_out
    (
      .clk                                         (video_clk),
      .lcd_data_format_adapter_1_out_data          (lcd_data_format_adapter_1_out_data),
      .lcd_data_format_adapter_1_out_empty         (lcd_data_format_adapter_1_out_empty),
      .lcd_data_format_adapter_1_out_endofpacket   (lcd_data_format_adapter_1_out_endofpacket),
      .lcd_data_format_adapter_1_out_ready         (lcd_data_format_adapter_1_out_ready),
      .lcd_data_format_adapter_1_out_startofpacket (lcd_data_format_adapter_1_out_startofpacket),
      .lcd_data_format_adapter_1_out_valid         (lcd_data_format_adapter_1_out_valid),
      .lcd_video_sequencer_in_ready_from_sa        (lcd_video_sequencer_in_ready_from_sa),
      .reset_n                                     (video_clk_reset_n)
    );

  lcd_data_format_adapter_1 the_lcd_data_format_adapter_1
    (
      .clk               (video_clk),
      .in_data           (lcd_data_format_adapter_1_in_data),
      .in_endofpacket    (lcd_data_format_adapter_1_in_endofpacket),
      .in_ready          (lcd_data_format_adapter_1_in_ready),
      .in_startofpacket  (lcd_data_format_adapter_1_in_startofpacket),
      .in_valid          (lcd_data_format_adapter_1_in_valid),
      .out_data          (lcd_data_format_adapter_1_out_data),
      .out_empty         (lcd_data_format_adapter_1_out_empty),
      .out_endofpacket   (lcd_data_format_adapter_1_out_endofpacket),
      .out_ready         (lcd_data_format_adapter_1_out_ready),
      .out_startofpacket (lcd_data_format_adapter_1_out_startofpacket),
      .out_valid         (lcd_data_format_adapter_1_out_valid),
      .reset_n           (lcd_data_format_adapter_1_in_reset_n)
    );

  lcd_i2c_cs_s1_arbitrator the_lcd_i2c_cs_s1
    (
      .clk                                                      (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1           (clock_crossing_bridge_m1_granted_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_latency_counter                 (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                   (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1 (clock_crossing_bridge_m1_qualified_request_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_read                            (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1   (clock_crossing_bridge_m1_read_data_valid_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1          (clock_crossing_bridge_m1_requests_lcd_i2c_cs_s1),
      .clock_crossing_bridge_m1_write                           (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                       (clock_crossing_bridge_m1_writedata),
      .d1_lcd_i2c_cs_s1_end_xfer                                (d1_lcd_i2c_cs_s1_end_xfer),
      .lcd_i2c_cs_s1_address                                    (lcd_i2c_cs_s1_address),
      .lcd_i2c_cs_s1_chipselect                                 (lcd_i2c_cs_s1_chipselect),
      .lcd_i2c_cs_s1_readdata                                   (lcd_i2c_cs_s1_readdata),
      .lcd_i2c_cs_s1_readdata_from_sa                           (lcd_i2c_cs_s1_readdata_from_sa),
      .lcd_i2c_cs_s1_reset_n                                    (lcd_i2c_cs_s1_reset_n),
      .lcd_i2c_cs_s1_write_n                                    (lcd_i2c_cs_s1_write_n),
      .lcd_i2c_cs_s1_writedata                                  (lcd_i2c_cs_s1_writedata),
      .reset_n                                                  (slow_clk_reset_n)
    );

  lcd_i2c_cs the_lcd_i2c_cs
    (
      .address    (lcd_i2c_cs_s1_address),
      .chipselect (lcd_i2c_cs_s1_chipselect),
      .clk        (slow_clk),
      .out_port   (out_port_from_the_lcd_i2c_cs),
      .readdata   (lcd_i2c_cs_s1_readdata),
      .reset_n    (lcd_i2c_cs_s1_reset_n),
      .write_n    (lcd_i2c_cs_s1_write_n),
      .writedata  (lcd_i2c_cs_s1_writedata)
    );

  lcd_i2c_dat_s1_arbitrator the_lcd_i2c_dat_s1
    (
      .clk                                                       (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                 (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1           (clock_crossing_bridge_m1_granted_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_latency_counter                  (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                    (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1 (clock_crossing_bridge_m1_qualified_request_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_read                             (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1   (clock_crossing_bridge_m1_read_data_valid_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1          (clock_crossing_bridge_m1_requests_lcd_i2c_dat_s1),
      .clock_crossing_bridge_m1_write                            (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                        (clock_crossing_bridge_m1_writedata),
      .d1_lcd_i2c_dat_s1_end_xfer                                (d1_lcd_i2c_dat_s1_end_xfer),
      .lcd_i2c_dat_s1_address                                    (lcd_i2c_dat_s1_address),
      .lcd_i2c_dat_s1_chipselect                                 (lcd_i2c_dat_s1_chipselect),
      .lcd_i2c_dat_s1_readdata                                   (lcd_i2c_dat_s1_readdata),
      .lcd_i2c_dat_s1_readdata_from_sa                           (lcd_i2c_dat_s1_readdata_from_sa),
      .lcd_i2c_dat_s1_reset_n                                    (lcd_i2c_dat_s1_reset_n),
      .lcd_i2c_dat_s1_write_n                                    (lcd_i2c_dat_s1_write_n),
      .lcd_i2c_dat_s1_writedata                                  (lcd_i2c_dat_s1_writedata),
      .reset_n                                                   (slow_clk_reset_n)
    );

  lcd_i2c_dat the_lcd_i2c_dat
    (
      .address    (lcd_i2c_dat_s1_address),
      .bidir_port (bidir_port_to_and_from_the_lcd_i2c_dat),
      .chipselect (lcd_i2c_dat_s1_chipselect),
      .clk        (slow_clk),
      .readdata   (lcd_i2c_dat_s1_readdata),
      .reset_n    (lcd_i2c_dat_s1_reset_n),
      .write_n    (lcd_i2c_dat_s1_write_n),
      .writedata  (lcd_i2c_dat_s1_writedata)
    );

  lcd_i2c_scl_s1_arbitrator the_lcd_i2c_scl_s1
    (
      .clk                                                       (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                 (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1           (clock_crossing_bridge_m1_granted_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_latency_counter                  (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                    (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1 (clock_crossing_bridge_m1_qualified_request_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_read                             (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1   (clock_crossing_bridge_m1_read_data_valid_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1          (clock_crossing_bridge_m1_requests_lcd_i2c_scl_s1),
      .clock_crossing_bridge_m1_write                            (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                        (clock_crossing_bridge_m1_writedata),
      .d1_lcd_i2c_scl_s1_end_xfer                                (d1_lcd_i2c_scl_s1_end_xfer),
      .lcd_i2c_scl_s1_address                                    (lcd_i2c_scl_s1_address),
      .lcd_i2c_scl_s1_chipselect                                 (lcd_i2c_scl_s1_chipselect),
      .lcd_i2c_scl_s1_readdata                                   (lcd_i2c_scl_s1_readdata),
      .lcd_i2c_scl_s1_readdata_from_sa                           (lcd_i2c_scl_s1_readdata_from_sa),
      .lcd_i2c_scl_s1_reset_n                                    (lcd_i2c_scl_s1_reset_n),
      .lcd_i2c_scl_s1_write_n                                    (lcd_i2c_scl_s1_write_n),
      .lcd_i2c_scl_s1_writedata                                  (lcd_i2c_scl_s1_writedata),
      .reset_n                                                   (slow_clk_reset_n)
    );

  lcd_i2c_scl the_lcd_i2c_scl
    (
      .address    (lcd_i2c_scl_s1_address),
      .chipselect (lcd_i2c_scl_s1_chipselect),
      .clk        (slow_clk),
      .out_port   (out_port_from_the_lcd_i2c_scl),
      .readdata   (lcd_i2c_scl_s1_readdata),
      .reset_n    (lcd_i2c_scl_s1_reset_n),
      .write_n    (lcd_i2c_scl_s1_write_n),
      .writedata  (lcd_i2c_scl_s1_writedata)
    );

  lcd_on_chip_memory_fifo_in_arbitrator the_lcd_on_chip_memory_fifo_in
    (
      .clk                                        (system_clk),
      .lcd_on_chip_memory_fifo_in_data            (lcd_on_chip_memory_fifo_in_data),
      .lcd_on_chip_memory_fifo_in_endofpacket     (lcd_on_chip_memory_fifo_in_endofpacket),
      .lcd_on_chip_memory_fifo_in_ready           (lcd_on_chip_memory_fifo_in_ready),
      .lcd_on_chip_memory_fifo_in_ready_from_sa   (lcd_on_chip_memory_fifo_in_ready_from_sa),
      .lcd_on_chip_memory_fifo_in_reset_n         (lcd_on_chip_memory_fifo_in_reset_n),
      .lcd_on_chip_memory_fifo_in_startofpacket   (lcd_on_chip_memory_fifo_in_startofpacket),
      .lcd_on_chip_memory_fifo_in_valid           (lcd_on_chip_memory_fifo_in_valid),
      .lcd_ta_formatter_to_fifo_out_data          (lcd_ta_formatter_to_fifo_out_data),
      .lcd_ta_formatter_to_fifo_out_endofpacket   (lcd_ta_formatter_to_fifo_out_endofpacket),
      .lcd_ta_formatter_to_fifo_out_startofpacket (lcd_ta_formatter_to_fifo_out_startofpacket),
      .lcd_ta_formatter_to_fifo_out_valid         (lcd_ta_formatter_to_fifo_out_valid),
      .reset_n                                    (system_clk_reset_n)
    );

  lcd_on_chip_memory_fifo_out_arbitrator the_lcd_on_chip_memory_fifo_out
    (
      .clk                                       (video_clk),
      .lcd_on_chip_memory_fifo_out_data          (lcd_on_chip_memory_fifo_out_data),
      .lcd_on_chip_memory_fifo_out_endofpacket   (lcd_on_chip_memory_fifo_out_endofpacket),
      .lcd_on_chip_memory_fifo_out_ready         (lcd_on_chip_memory_fifo_out_ready),
      .lcd_on_chip_memory_fifo_out_reset_n       (lcd_on_chip_memory_fifo_out_reset_n),
      .lcd_on_chip_memory_fifo_out_startofpacket (lcd_on_chip_memory_fifo_out_startofpacket),
      .lcd_on_chip_memory_fifo_out_valid         (lcd_on_chip_memory_fifo_out_valid),
      .lcd_ta_fifo_to_sequencer_in_ready_from_sa (lcd_ta_fifo_to_sequencer_in_ready_from_sa),
      .reset_n                                   (video_clk_reset_n)
    );

  lcd_on_chip_memory_fifo the_lcd_on_chip_memory_fifo
    (
      .avalonst_sink_data            (lcd_on_chip_memory_fifo_in_data),
      .avalonst_sink_endofpacket     (lcd_on_chip_memory_fifo_in_endofpacket),
      .avalonst_sink_ready           (lcd_on_chip_memory_fifo_in_ready),
      .avalonst_sink_startofpacket   (lcd_on_chip_memory_fifo_in_startofpacket),
      .avalonst_sink_valid           (lcd_on_chip_memory_fifo_in_valid),
      .avalonst_source_data          (lcd_on_chip_memory_fifo_out_data),
      .avalonst_source_endofpacket   (lcd_on_chip_memory_fifo_out_endofpacket),
      .avalonst_source_ready         (lcd_on_chip_memory_fifo_out_ready),
      .avalonst_source_startofpacket (lcd_on_chip_memory_fifo_out_startofpacket),
      .avalonst_source_valid         (lcd_on_chip_memory_fifo_out_valid),
      .rdclock                       (video_clk),
      .rdreset_n                     (lcd_on_chip_memory_fifo_out_reset_n),
      .wrclock                       (system_clk),
      .wrreset_n                     (lcd_on_chip_memory_fifo_in_reset_n)
    );

  lcd_pixel_converter_in_arbitrator the_lcd_pixel_converter_in
    (
      .clk                                  (system_clk),
      .lcd_pixel_converter_in_data          (lcd_pixel_converter_in_data),
      .lcd_pixel_converter_in_empty         (lcd_pixel_converter_in_empty),
      .lcd_pixel_converter_in_endofpacket   (lcd_pixel_converter_in_endofpacket),
      .lcd_pixel_converter_in_ready         (lcd_pixel_converter_in_ready),
      .lcd_pixel_converter_in_ready_from_sa (lcd_pixel_converter_in_ready_from_sa),
      .lcd_pixel_converter_in_reset_n       (lcd_pixel_converter_in_reset_n),
      .lcd_pixel_converter_in_startofpacket (lcd_pixel_converter_in_startofpacket),
      .lcd_pixel_converter_in_valid         (lcd_pixel_converter_in_valid),
      .lcd_sgdma_out_data                   (lcd_sgdma_out_data),
      .lcd_sgdma_out_empty                  (lcd_sgdma_out_empty),
      .lcd_sgdma_out_endofpacket            (lcd_sgdma_out_endofpacket),
      .lcd_sgdma_out_startofpacket          (lcd_sgdma_out_startofpacket),
      .lcd_sgdma_out_valid                  (lcd_sgdma_out_valid),
      .reset_n                              (system_clk_reset_n)
    );

  lcd_pixel_converter_out_arbitrator the_lcd_pixel_converter_out
    (
      .clk                                      (system_clk),
      .lcd_data_format_adapter_in_ready_from_sa (lcd_data_format_adapter_in_ready_from_sa),
      .lcd_pixel_converter_out_data             (lcd_pixel_converter_out_data),
      .lcd_pixel_converter_out_empty            (lcd_pixel_converter_out_empty),
      .lcd_pixel_converter_out_endofpacket      (lcd_pixel_converter_out_endofpacket),
      .lcd_pixel_converter_out_ready            (lcd_pixel_converter_out_ready),
      .lcd_pixel_converter_out_startofpacket    (lcd_pixel_converter_out_startofpacket),
      .lcd_pixel_converter_out_valid            (lcd_pixel_converter_out_valid),
      .reset_n                                  (system_clk_reset_n)
    );

  lcd_pixel_converter the_lcd_pixel_converter
    (
      .clk       (system_clk),
      .data_in   (lcd_pixel_converter_in_data),
      .data_out  (lcd_pixel_converter_out_data),
      .empty_in  (lcd_pixel_converter_in_empty),
      .empty_out (lcd_pixel_converter_out_empty),
      .eop_in    (lcd_pixel_converter_in_endofpacket),
      .eop_out   (lcd_pixel_converter_out_endofpacket),
      .ready_in  (lcd_pixel_converter_out_ready),
      .ready_out (lcd_pixel_converter_in_ready),
      .reset_n   (lcd_pixel_converter_in_reset_n),
      .sop_in    (lcd_pixel_converter_in_startofpacket),
      .sop_out   (lcd_pixel_converter_out_startofpacket),
      .valid_in  (lcd_pixel_converter_in_valid),
      .valid_out (lcd_pixel_converter_out_valid)
    );

  lcd_sgdma_csr_arbitrator the_lcd_sgdma_csr
    (
      .clk                                                                               (system_clk),
      .d1_lcd_sgdma_csr_end_xfer                                                         (d1_lcd_sgdma_csr_end_xfer),
      .lcd_sgdma_csr_address                                                             (lcd_sgdma_csr_address),
      .lcd_sgdma_csr_chipselect                                                          (lcd_sgdma_csr_chipselect),
      .lcd_sgdma_csr_irq                                                                 (lcd_sgdma_csr_irq),
      .lcd_sgdma_csr_irq_from_sa                                                         (lcd_sgdma_csr_irq_from_sa),
      .lcd_sgdma_csr_read                                                                (lcd_sgdma_csr_read),
      .lcd_sgdma_csr_readdata                                                            (lcd_sgdma_csr_readdata),
      .lcd_sgdma_csr_readdata_from_sa                                                    (lcd_sgdma_csr_readdata_from_sa),
      .lcd_sgdma_csr_reset_n                                                             (lcd_sgdma_csr_reset_n),
      .lcd_sgdma_csr_write                                                               (lcd_sgdma_csr_write),
      .lcd_sgdma_csr_writedata                                                           (lcd_sgdma_csr_writedata),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_lcd_sgdma_csr                                          (pipeline_bridge_m1_granted_lcd_sgdma_csr),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_lcd_sgdma_csr                                (pipeline_bridge_m1_qualified_request_lcd_sgdma_csr),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr                                  (pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr),
      .pipeline_bridge_m1_requests_lcd_sgdma_csr                                         (pipeline_bridge_m1_requests_lcd_sgdma_csr),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  lcd_sgdma_descriptor_read_arbitrator the_lcd_sgdma_descriptor_read
    (
      .clk                                                              (system_clk),
      .d1_descriptor_memory_s2_end_xfer                                 (d1_descriptor_memory_s2_end_xfer),
      .descriptor_memory_s2_readdata_from_sa                            (descriptor_memory_s2_readdata_from_sa),
      .lcd_sgdma_descriptor_read_address                                (lcd_sgdma_descriptor_read_address),
      .lcd_sgdma_descriptor_read_address_to_slave                       (lcd_sgdma_descriptor_read_address_to_slave),
      .lcd_sgdma_descriptor_read_granted_descriptor_memory_s2           (lcd_sgdma_descriptor_read_granted_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_latency_counter                        (lcd_sgdma_descriptor_read_latency_counter),
      .lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2 (lcd_sgdma_descriptor_read_qualified_request_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_read                                   (lcd_sgdma_descriptor_read_read),
      .lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2   (lcd_sgdma_descriptor_read_read_data_valid_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_readdata                               (lcd_sgdma_descriptor_read_readdata),
      .lcd_sgdma_descriptor_read_readdatavalid                          (lcd_sgdma_descriptor_read_readdatavalid),
      .lcd_sgdma_descriptor_read_requests_descriptor_memory_s2          (lcd_sgdma_descriptor_read_requests_descriptor_memory_s2),
      .lcd_sgdma_descriptor_read_waitrequest                            (lcd_sgdma_descriptor_read_waitrequest),
      .reset_n                                                          (system_clk_reset_n)
    );

  lcd_sgdma_descriptor_write_arbitrator the_lcd_sgdma_descriptor_write
    (
      .clk                                                               (system_clk),
      .d1_descriptor_memory_s2_end_xfer                                  (d1_descriptor_memory_s2_end_xfer),
      .lcd_sgdma_descriptor_write_address                                (lcd_sgdma_descriptor_write_address),
      .lcd_sgdma_descriptor_write_address_to_slave                       (lcd_sgdma_descriptor_write_address_to_slave),
      .lcd_sgdma_descriptor_write_granted_descriptor_memory_s2           (lcd_sgdma_descriptor_write_granted_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2 (lcd_sgdma_descriptor_write_qualified_request_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_requests_descriptor_memory_s2          (lcd_sgdma_descriptor_write_requests_descriptor_memory_s2),
      .lcd_sgdma_descriptor_write_waitrequest                            (lcd_sgdma_descriptor_write_waitrequest),
      .lcd_sgdma_descriptor_write_write                                  (lcd_sgdma_descriptor_write_write),
      .lcd_sgdma_descriptor_write_writedata                              (lcd_sgdma_descriptor_write_writedata),
      .reset_n                                                           (system_clk_reset_n)
    );

  lcd_sgdma_m_read_arbitrator the_lcd_sgdma_m_read
    (
      .clk                                                                             (system_clk),
      .d1_frame_buffer_pipeline_bridge_s1_end_xfer                                     (d1_frame_buffer_pipeline_bridge_s1_end_xfer),
      .frame_buffer_pipeline_bridge_s1_readdata_from_sa                                (frame_buffer_pipeline_bridge_s1_readdata_from_sa),
      .frame_buffer_pipeline_bridge_s1_waitrequest_from_sa                             (frame_buffer_pipeline_bridge_s1_waitrequest_from_sa),
      .lcd_sgdma_m_read_address                                                        (lcd_sgdma_m_read_address),
      .lcd_sgdma_m_read_address_to_slave                                               (lcd_sgdma_m_read_address_to_slave),
      .lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1                        (lcd_sgdma_m_read_granted_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_latency_counter                                                (lcd_sgdma_m_read_latency_counter),
      .lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1              (lcd_sgdma_m_read_qualified_request_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_read                                                           (lcd_sgdma_m_read_read),
      .lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1                (lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (lcd_sgdma_m_read_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .lcd_sgdma_m_read_readdata                                                       (lcd_sgdma_m_read_readdata),
      .lcd_sgdma_m_read_readdatavalid                                                  (lcd_sgdma_m_read_readdatavalid),
      .lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1                       (lcd_sgdma_m_read_requests_frame_buffer_pipeline_bridge_s1),
      .lcd_sgdma_m_read_waitrequest                                                    (lcd_sgdma_m_read_waitrequest),
      .reset_n                                                                         (system_clk_reset_n)
    );

  lcd_sgdma_out_arbitrator the_lcd_sgdma_out
    (
      .clk                                  (system_clk),
      .lcd_pixel_converter_in_ready_from_sa (lcd_pixel_converter_in_ready_from_sa),
      .lcd_sgdma_out_data                   (lcd_sgdma_out_data),
      .lcd_sgdma_out_empty                  (lcd_sgdma_out_empty),
      .lcd_sgdma_out_endofpacket            (lcd_sgdma_out_endofpacket),
      .lcd_sgdma_out_ready                  (lcd_sgdma_out_ready),
      .lcd_sgdma_out_startofpacket          (lcd_sgdma_out_startofpacket),
      .lcd_sgdma_out_valid                  (lcd_sgdma_out_valid),
      .reset_n                              (system_clk_reset_n)
    );

  lcd_sgdma the_lcd_sgdma
    (
      .clk                           (system_clk),
      .csr_address                   (lcd_sgdma_csr_address),
      .csr_chipselect                (lcd_sgdma_csr_chipselect),
      .csr_irq                       (lcd_sgdma_csr_irq),
      .csr_read                      (lcd_sgdma_csr_read),
      .csr_readdata                  (lcd_sgdma_csr_readdata),
      .csr_write                     (lcd_sgdma_csr_write),
      .csr_writedata                 (lcd_sgdma_csr_writedata),
      .descriptor_read_address       (lcd_sgdma_descriptor_read_address),
      .descriptor_read_read          (lcd_sgdma_descriptor_read_read),
      .descriptor_read_readdata      (lcd_sgdma_descriptor_read_readdata),
      .descriptor_read_readdatavalid (lcd_sgdma_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (lcd_sgdma_descriptor_read_waitrequest),
      .descriptor_write_address      (lcd_sgdma_descriptor_write_address),
      .descriptor_write_waitrequest  (lcd_sgdma_descriptor_write_waitrequest),
      .descriptor_write_write        (lcd_sgdma_descriptor_write_write),
      .descriptor_write_writedata    (lcd_sgdma_descriptor_write_writedata),
      .m_read_address                (lcd_sgdma_m_read_address),
      .m_read_read                   (lcd_sgdma_m_read_read),
      .m_read_readdata               (lcd_sgdma_m_read_readdata),
      .m_read_readdatavalid          (lcd_sgdma_m_read_readdatavalid),
      .m_read_waitrequest            (lcd_sgdma_m_read_waitrequest),
      .out_data                      (lcd_sgdma_out_data),
      .out_empty                     (lcd_sgdma_out_empty),
      .out_endofpacket               (lcd_sgdma_out_endofpacket),
      .out_ready                     (lcd_sgdma_out_ready),
      .out_startofpacket             (lcd_sgdma_out_startofpacket),
      .out_valid                     (lcd_sgdma_out_valid),
      .system_reset_n                (lcd_sgdma_csr_reset_n)
    );

  lcd_ta_fifo_to_sequencer_in_arbitrator the_lcd_ta_fifo_to_sequencer_in
    (
      .clk                                       (video_clk),
      .lcd_on_chip_memory_fifo_out_data          (lcd_on_chip_memory_fifo_out_data),
      .lcd_on_chip_memory_fifo_out_endofpacket   (lcd_on_chip_memory_fifo_out_endofpacket),
      .lcd_on_chip_memory_fifo_out_startofpacket (lcd_on_chip_memory_fifo_out_startofpacket),
      .lcd_on_chip_memory_fifo_out_valid         (lcd_on_chip_memory_fifo_out_valid),
      .lcd_ta_fifo_to_sequencer_in_data          (lcd_ta_fifo_to_sequencer_in_data),
      .lcd_ta_fifo_to_sequencer_in_endofpacket   (lcd_ta_fifo_to_sequencer_in_endofpacket),
      .lcd_ta_fifo_to_sequencer_in_ready         (lcd_ta_fifo_to_sequencer_in_ready),
      .lcd_ta_fifo_to_sequencer_in_ready_from_sa (lcd_ta_fifo_to_sequencer_in_ready_from_sa),
      .lcd_ta_fifo_to_sequencer_in_reset_n       (lcd_ta_fifo_to_sequencer_in_reset_n),
      .lcd_ta_fifo_to_sequencer_in_startofpacket (lcd_ta_fifo_to_sequencer_in_startofpacket),
      .lcd_ta_fifo_to_sequencer_in_valid         (lcd_ta_fifo_to_sequencer_in_valid),
      .reset_n                                   (video_clk_reset_n)
    );

  lcd_ta_fifo_to_sequencer_out_arbitrator the_lcd_ta_fifo_to_sequencer_out
    (
      .clk                                        (video_clk),
      .lcd_data_format_adapter_1_in_ready_from_sa (lcd_data_format_adapter_1_in_ready_from_sa),
      .lcd_ta_fifo_to_sequencer_out_data          (lcd_ta_fifo_to_sequencer_out_data),
      .lcd_ta_fifo_to_sequencer_out_endofpacket   (lcd_ta_fifo_to_sequencer_out_endofpacket),
      .lcd_ta_fifo_to_sequencer_out_ready         (lcd_ta_fifo_to_sequencer_out_ready),
      .lcd_ta_fifo_to_sequencer_out_startofpacket (lcd_ta_fifo_to_sequencer_out_startofpacket),
      .lcd_ta_fifo_to_sequencer_out_valid         (lcd_ta_fifo_to_sequencer_out_valid),
      .reset_n                                    (video_clk_reset_n)
    );

  lcd_ta_fifo_to_sequencer the_lcd_ta_fifo_to_sequencer
    (
      .clk               (video_clk),
      .in_data           (lcd_ta_fifo_to_sequencer_in_data),
      .in_endofpacket    (lcd_ta_fifo_to_sequencer_in_endofpacket),
      .in_ready          (lcd_ta_fifo_to_sequencer_in_ready),
      .in_startofpacket  (lcd_ta_fifo_to_sequencer_in_startofpacket),
      .in_valid          (lcd_ta_fifo_to_sequencer_in_valid),
      .out_data          (lcd_ta_fifo_to_sequencer_out_data),
      .out_endofpacket   (lcd_ta_fifo_to_sequencer_out_endofpacket),
      .out_ready         (lcd_ta_fifo_to_sequencer_out_ready),
      .out_startofpacket (lcd_ta_fifo_to_sequencer_out_startofpacket),
      .out_valid         (lcd_ta_fifo_to_sequencer_out_valid),
      .reset_n           (lcd_ta_fifo_to_sequencer_in_reset_n)
    );

  lcd_ta_formatter_to_fifo_in_arbitrator the_lcd_ta_formatter_to_fifo_in
    (
      .clk                                       (system_clk),
      .lcd_data_format_adapter_out_data          (lcd_data_format_adapter_out_data),
      .lcd_data_format_adapter_out_endofpacket   (lcd_data_format_adapter_out_endofpacket),
      .lcd_data_format_adapter_out_startofpacket (lcd_data_format_adapter_out_startofpacket),
      .lcd_data_format_adapter_out_valid         (lcd_data_format_adapter_out_valid),
      .lcd_ta_formatter_to_fifo_in_data          (lcd_ta_formatter_to_fifo_in_data),
      .lcd_ta_formatter_to_fifo_in_endofpacket   (lcd_ta_formatter_to_fifo_in_endofpacket),
      .lcd_ta_formatter_to_fifo_in_ready         (lcd_ta_formatter_to_fifo_in_ready),
      .lcd_ta_formatter_to_fifo_in_ready_from_sa (lcd_ta_formatter_to_fifo_in_ready_from_sa),
      .lcd_ta_formatter_to_fifo_in_reset_n       (lcd_ta_formatter_to_fifo_in_reset_n),
      .lcd_ta_formatter_to_fifo_in_startofpacket (lcd_ta_formatter_to_fifo_in_startofpacket),
      .lcd_ta_formatter_to_fifo_in_valid         (lcd_ta_formatter_to_fifo_in_valid),
      .reset_n                                   (system_clk_reset_n)
    );

  lcd_ta_formatter_to_fifo_out_arbitrator the_lcd_ta_formatter_to_fifo_out
    (
      .clk                                        (system_clk),
      .lcd_on_chip_memory_fifo_in_ready_from_sa   (lcd_on_chip_memory_fifo_in_ready_from_sa),
      .lcd_ta_formatter_to_fifo_out_data          (lcd_ta_formatter_to_fifo_out_data),
      .lcd_ta_formatter_to_fifo_out_endofpacket   (lcd_ta_formatter_to_fifo_out_endofpacket),
      .lcd_ta_formatter_to_fifo_out_ready         (lcd_ta_formatter_to_fifo_out_ready),
      .lcd_ta_formatter_to_fifo_out_startofpacket (lcd_ta_formatter_to_fifo_out_startofpacket),
      .lcd_ta_formatter_to_fifo_out_valid         (lcd_ta_formatter_to_fifo_out_valid),
      .reset_n                                    (system_clk_reset_n)
    );

  lcd_ta_formatter_to_fifo the_lcd_ta_formatter_to_fifo
    (
      .clk               (system_clk),
      .in_data           (lcd_ta_formatter_to_fifo_in_data),
      .in_endofpacket    (lcd_ta_formatter_to_fifo_in_endofpacket),
      .in_ready          (lcd_ta_formatter_to_fifo_in_ready),
      .in_startofpacket  (lcd_ta_formatter_to_fifo_in_startofpacket),
      .in_valid          (lcd_ta_formatter_to_fifo_in_valid),
      .out_data          (lcd_ta_formatter_to_fifo_out_data),
      .out_endofpacket   (lcd_ta_formatter_to_fifo_out_endofpacket),
      .out_ready         (lcd_ta_formatter_to_fifo_out_ready),
      .out_startofpacket (lcd_ta_formatter_to_fifo_out_startofpacket),
      .out_valid         (lcd_ta_formatter_to_fifo_out_valid),
      .reset_n           (lcd_ta_formatter_to_fifo_in_reset_n)
    );

  lcd_video_sequencer_in_arbitrator the_lcd_video_sequencer_in
    (
      .clk                                         (video_clk),
      .lcd_data_format_adapter_1_out_data          (lcd_data_format_adapter_1_out_data),
      .lcd_data_format_adapter_1_out_empty         (lcd_data_format_adapter_1_out_empty),
      .lcd_data_format_adapter_1_out_endofpacket   (lcd_data_format_adapter_1_out_endofpacket),
      .lcd_data_format_adapter_1_out_startofpacket (lcd_data_format_adapter_1_out_startofpacket),
      .lcd_data_format_adapter_1_out_valid         (lcd_data_format_adapter_1_out_valid),
      .lcd_video_sequencer_in_data                 (lcd_video_sequencer_in_data),
      .lcd_video_sequencer_in_empty                (lcd_video_sequencer_in_empty),
      .lcd_video_sequencer_in_endofpacket          (lcd_video_sequencer_in_endofpacket),
      .lcd_video_sequencer_in_ready                (lcd_video_sequencer_in_ready),
      .lcd_video_sequencer_in_ready_from_sa        (lcd_video_sequencer_in_ready_from_sa),
      .lcd_video_sequencer_in_reset_n              (lcd_video_sequencer_in_reset_n),
      .lcd_video_sequencer_in_startofpacket        (lcd_video_sequencer_in_startofpacket),
      .lcd_video_sequencer_in_valid                (lcd_video_sequencer_in_valid),
      .reset_n                                     (video_clk_reset_n)
    );

  lcd_video_sequencer the_lcd_video_sequencer
    (
      .DEN     (DEN_from_the_lcd_video_sequencer),
      .HD      (HD_from_the_lcd_video_sequencer),
      .RGB_OUT (RGB_OUT_from_the_lcd_video_sequencer),
      .VD      (VD_from_the_lcd_video_sequencer),
      .clk     (video_clk),
      .data    (lcd_video_sequencer_in_data),
      .empty   (lcd_video_sequencer_in_empty),
      .eop     (lcd_video_sequencer_in_endofpacket),
      .ready   (lcd_video_sequencer_in_ready),
      .reset_n (lcd_video_sequencer_in_reset_n),
      .sop     (lcd_video_sequencer_in_startofpacket),
      .valid   (lcd_video_sequencer_in_valid)
    );

  pio_id_eeprom_dat_s1_arbitrator the_pio_id_eeprom_dat_s1
    (
      .clk                                                             (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                       (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1           (clock_crossing_bridge_m1_granted_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_latency_counter                        (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                          (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1 (clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_read                                   (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1   (clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1          (clock_crossing_bridge_m1_requests_pio_id_eeprom_dat_s1),
      .clock_crossing_bridge_m1_write                                  (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                              (clock_crossing_bridge_m1_writedata),
      .d1_pio_id_eeprom_dat_s1_end_xfer                                (d1_pio_id_eeprom_dat_s1_end_xfer),
      .pio_id_eeprom_dat_s1_address                                    (pio_id_eeprom_dat_s1_address),
      .pio_id_eeprom_dat_s1_chipselect                                 (pio_id_eeprom_dat_s1_chipselect),
      .pio_id_eeprom_dat_s1_readdata                                   (pio_id_eeprom_dat_s1_readdata),
      .pio_id_eeprom_dat_s1_readdata_from_sa                           (pio_id_eeprom_dat_s1_readdata_from_sa),
      .pio_id_eeprom_dat_s1_reset_n                                    (pio_id_eeprom_dat_s1_reset_n),
      .pio_id_eeprom_dat_s1_write_n                                    (pio_id_eeprom_dat_s1_write_n),
      .pio_id_eeprom_dat_s1_writedata                                  (pio_id_eeprom_dat_s1_writedata),
      .reset_n                                                         (slow_clk_reset_n)
    );

  pio_id_eeprom_dat the_pio_id_eeprom_dat
    (
      .address    (pio_id_eeprom_dat_s1_address),
      .bidir_port (bidir_port_to_and_from_the_pio_id_eeprom_dat),
      .chipselect (pio_id_eeprom_dat_s1_chipselect),
      .clk        (slow_clk),
      .readdata   (pio_id_eeprom_dat_s1_readdata),
      .reset_n    (pio_id_eeprom_dat_s1_reset_n),
      .write_n    (pio_id_eeprom_dat_s1_write_n),
      .writedata  (pio_id_eeprom_dat_s1_writedata)
    );

  pio_id_eeprom_scl_s1_arbitrator the_pio_id_eeprom_scl_s1
    (
      .clk                                                             (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                       (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1           (clock_crossing_bridge_m1_granted_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_latency_counter                        (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                          (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1 (clock_crossing_bridge_m1_qualified_request_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_read                                   (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1   (clock_crossing_bridge_m1_read_data_valid_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1          (clock_crossing_bridge_m1_requests_pio_id_eeprom_scl_s1),
      .clock_crossing_bridge_m1_write                                  (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                              (clock_crossing_bridge_m1_writedata),
      .d1_pio_id_eeprom_scl_s1_end_xfer                                (d1_pio_id_eeprom_scl_s1_end_xfer),
      .pio_id_eeprom_scl_s1_address                                    (pio_id_eeprom_scl_s1_address),
      .pio_id_eeprom_scl_s1_chipselect                                 (pio_id_eeprom_scl_s1_chipselect),
      .pio_id_eeprom_scl_s1_readdata                                   (pio_id_eeprom_scl_s1_readdata),
      .pio_id_eeprom_scl_s1_readdata_from_sa                           (pio_id_eeprom_scl_s1_readdata_from_sa),
      .pio_id_eeprom_scl_s1_reset_n                                    (pio_id_eeprom_scl_s1_reset_n),
      .pio_id_eeprom_scl_s1_write_n                                    (pio_id_eeprom_scl_s1_write_n),
      .pio_id_eeprom_scl_s1_writedata                                  (pio_id_eeprom_scl_s1_writedata),
      .reset_n                                                         (slow_clk_reset_n)
    );

  pio_id_eeprom_scl the_pio_id_eeprom_scl
    (
      .address    (pio_id_eeprom_scl_s1_address),
      .chipselect (pio_id_eeprom_scl_s1_chipselect),
      .clk        (slow_clk),
      .out_port   (out_port_from_the_pio_id_eeprom_scl),
      .readdata   (pio_id_eeprom_scl_s1_readdata),
      .reset_n    (pio_id_eeprom_scl_s1_reset_n),
      .write_n    (pio_id_eeprom_scl_s1_write_n),
      .writedata  (pio_id_eeprom_scl_s1_writedata)
    );

  pipeline_bridge_s1_arbitrator the_pipeline_bridge_s1
    (
      .clk                                                                      (system_clk),
      .cpu_data_master_address_to_slave                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                               (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                              (cpu_data_master_debugaccess),
      .cpu_data_master_granted_pipeline_bridge_s1                               (cpu_data_master_granted_pipeline_bridge_s1),
      .cpu_data_master_latency_counter                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_pipeline_bridge_s1                     (cpu_data_master_qualified_request_pipeline_bridge_s1),
      .cpu_data_master_read                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_pipeline_bridge_s1                       (cpu_data_master_read_data_valid_pipeline_bridge_s1),
      .cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register        (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register),
      .cpu_data_master_requests_pipeline_bridge_s1                              (cpu_data_master_requests_pipeline_bridge_s1),
      .cpu_data_master_write                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                  (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_pipeline_bridge_s1                        (cpu_instruction_master_granted_pipeline_bridge_s1),
      .cpu_instruction_master_latency_counter                                   (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_pipeline_bridge_s1              (cpu_instruction_master_qualified_request_pipeline_bridge_s1),
      .cpu_instruction_master_read                                              (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_s1                (cpu_instruction_master_read_data_valid_pipeline_bridge_s1),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register (cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register),
      .cpu_instruction_master_requests_pipeline_bridge_s1                       (cpu_instruction_master_requests_pipeline_bridge_s1),
      .d1_pipeline_bridge_s1_end_xfer                                           (d1_pipeline_bridge_s1_end_xfer),
      .pipeline_bridge_s1_address                                               (pipeline_bridge_s1_address),
      .pipeline_bridge_s1_arbiterlock                                           (pipeline_bridge_s1_arbiterlock),
      .pipeline_bridge_s1_arbiterlock2                                          (pipeline_bridge_s1_arbiterlock2),
      .pipeline_bridge_s1_burstcount                                            (pipeline_bridge_s1_burstcount),
      .pipeline_bridge_s1_byteenable                                            (pipeline_bridge_s1_byteenable),
      .pipeline_bridge_s1_chipselect                                            (pipeline_bridge_s1_chipselect),
      .pipeline_bridge_s1_debugaccess                                           (pipeline_bridge_s1_debugaccess),
      .pipeline_bridge_s1_endofpacket                                           (pipeline_bridge_s1_endofpacket),
      .pipeline_bridge_s1_endofpacket_from_sa                                   (pipeline_bridge_s1_endofpacket_from_sa),
      .pipeline_bridge_s1_nativeaddress                                         (pipeline_bridge_s1_nativeaddress),
      .pipeline_bridge_s1_read                                                  (pipeline_bridge_s1_read),
      .pipeline_bridge_s1_readdata                                              (pipeline_bridge_s1_readdata),
      .pipeline_bridge_s1_readdata_from_sa                                      (pipeline_bridge_s1_readdata_from_sa),
      .pipeline_bridge_s1_readdatavalid                                         (pipeline_bridge_s1_readdatavalid),
      .pipeline_bridge_s1_reset_n                                               (pipeline_bridge_s1_reset_n),
      .pipeline_bridge_s1_waitrequest                                           (pipeline_bridge_s1_waitrequest),
      .pipeline_bridge_s1_waitrequest_from_sa                                   (pipeline_bridge_s1_waitrequest_from_sa),
      .pipeline_bridge_s1_write                                                 (pipeline_bridge_s1_write),
      .pipeline_bridge_s1_writedata                                             (pipeline_bridge_s1_writedata),
      .reset_n                                                                  (system_clk_reset_n)
    );

  pipeline_bridge_m1_arbitrator the_pipeline_bridge_m1
    (
      .clk                                                                               (system_clk),
      .clock_crossing_bridge_s1_endofpacket_from_sa                                      (clock_crossing_bridge_s1_endofpacket_from_sa),
      .clock_crossing_bridge_s1_readdata_from_sa                                         (clock_crossing_bridge_s1_readdata_from_sa),
      .clock_crossing_bridge_s1_waitrequest_from_sa                                      (clock_crossing_bridge_s1_waitrequest_from_sa),
      .colour_lookup_table_s1_readdata_from_sa                                           (colour_lookup_table_s1_readdata_from_sa),
      .cpu_jtag_debug_module_readdata_from_sa                                            (cpu_jtag_debug_module_readdata_from_sa),
      .d1_clock_crossing_bridge_s1_end_xfer                                              (d1_clock_crossing_bridge_s1_end_xfer),
      .d1_colour_lookup_table_s1_end_xfer                                                (d1_colour_lookup_table_s1_end_xfer),
      .d1_cpu_jtag_debug_module_end_xfer                                                 (d1_cpu_jtag_debug_module_end_xfer),
      .d1_descriptor_memory_s1_end_xfer                                                  (d1_descriptor_memory_s1_end_xfer),
      .d1_flash_ssram_pipeline_bridge_s1_end_xfer                                        (d1_flash_ssram_pipeline_bridge_s1_end_xfer),
      .d1_frame_buffer_pipeline_bridge_s1_end_xfer                                       (d1_frame_buffer_pipeline_bridge_s1_end_xfer),
      .d1_lcd_sgdma_csr_end_xfer                                                         (d1_lcd_sgdma_csr_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                                             (descriptor_memory_s1_readdata_from_sa),
      .flash_ssram_pipeline_bridge_s1_endofpacket_from_sa                                (flash_ssram_pipeline_bridge_s1_endofpacket_from_sa),
      .flash_ssram_pipeline_bridge_s1_readdata_from_sa                                   (flash_ssram_pipeline_bridge_s1_readdata_from_sa),
      .flash_ssram_pipeline_bridge_s1_waitrequest_from_sa                                (flash_ssram_pipeline_bridge_s1_waitrequest_from_sa),
      .frame_buffer_pipeline_bridge_s1_endofpacket_from_sa                               (frame_buffer_pipeline_bridge_s1_endofpacket_from_sa),
      .frame_buffer_pipeline_bridge_s1_readdata_from_sa                                  (frame_buffer_pipeline_bridge_s1_readdata_from_sa),
      .frame_buffer_pipeline_bridge_s1_waitrequest_from_sa                               (frame_buffer_pipeline_bridge_s1_waitrequest_from_sa),
      .lcd_sgdma_csr_readdata_from_sa                                                    (lcd_sgdma_csr_readdata_from_sa),
      .pipeline_bridge_m1_address                                                        (pipeline_bridge_m1_address),
      .pipeline_bridge_m1_address_to_slave                                               (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                                     (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                                     (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                                     (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_endofpacket                                                    (pipeline_bridge_m1_endofpacket),
      .pipeline_bridge_m1_granted_clock_crossing_bridge_s1                               (pipeline_bridge_m1_granted_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_granted_colour_lookup_table_s1                                 (pipeline_bridge_m1_granted_colour_lookup_table_s1),
      .pipeline_bridge_m1_granted_cpu_jtag_debug_module                                  (pipeline_bridge_m1_granted_cpu_jtag_debug_module),
      .pipeline_bridge_m1_granted_descriptor_memory_s1                                   (pipeline_bridge_m1_granted_descriptor_memory_s1),
      .pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1                         (pipeline_bridge_m1_granted_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1                        (pipeline_bridge_m1_granted_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_granted_lcd_sgdma_csr                                          (pipeline_bridge_m1_granted_lcd_sgdma_csr),
      .pipeline_bridge_m1_latency_counter                                                (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1                     (pipeline_bridge_m1_qualified_request_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_qualified_request_colour_lookup_table_s1                       (pipeline_bridge_m1_qualified_request_colour_lookup_table_s1),
      .pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module                        (pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module),
      .pipeline_bridge_m1_qualified_request_descriptor_memory_s1                         (pipeline_bridge_m1_qualified_request_descriptor_memory_s1),
      .pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1               (pipeline_bridge_m1_qualified_request_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1              (pipeline_bridge_m1_qualified_request_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_qualified_request_lcd_sgdma_csr                                (pipeline_bridge_m1_qualified_request_lcd_sgdma_csr),
      .pipeline_bridge_m1_read                                                           (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1                       (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register        (pipeline_bridge_m1_read_data_valid_clock_crossing_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1                         (pipeline_bridge_m1_read_data_valid_colour_lookup_table_s1),
      .pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module                          (pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module),
      .pipeline_bridge_m1_read_data_valid_descriptor_memory_s1                           (pipeline_bridge_m1_read_data_valid_descriptor_memory_s1),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1                 (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register  (pipeline_bridge_m1_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1                (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register (pipeline_bridge_m1_read_data_valid_frame_buffer_pipeline_bridge_s1_shift_register),
      .pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr                                  (pipeline_bridge_m1_read_data_valid_lcd_sgdma_csr),
      .pipeline_bridge_m1_readdata                                                       (pipeline_bridge_m1_readdata),
      .pipeline_bridge_m1_readdatavalid                                                  (pipeline_bridge_m1_readdatavalid),
      .pipeline_bridge_m1_requests_clock_crossing_bridge_s1                              (pipeline_bridge_m1_requests_clock_crossing_bridge_s1),
      .pipeline_bridge_m1_requests_colour_lookup_table_s1                                (pipeline_bridge_m1_requests_colour_lookup_table_s1),
      .pipeline_bridge_m1_requests_cpu_jtag_debug_module                                 (pipeline_bridge_m1_requests_cpu_jtag_debug_module),
      .pipeline_bridge_m1_requests_descriptor_memory_s1                                  (pipeline_bridge_m1_requests_descriptor_memory_s1),
      .pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1                        (pipeline_bridge_m1_requests_flash_ssram_pipeline_bridge_s1),
      .pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1                       (pipeline_bridge_m1_requests_frame_buffer_pipeline_bridge_s1),
      .pipeline_bridge_m1_requests_lcd_sgdma_csr                                         (pipeline_bridge_m1_requests_lcd_sgdma_csr),
      .pipeline_bridge_m1_waitrequest                                                    (pipeline_bridge_m1_waitrequest),
      .pipeline_bridge_m1_write                                                          (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                                      (pipeline_bridge_m1_writedata),
      .reset_n                                                                           (system_clk_reset_n)
    );

  pipeline_bridge the_pipeline_bridge
    (
      .clk              (system_clk),
      .m1_address       (pipeline_bridge_m1_address),
      .m1_burstcount    (pipeline_bridge_m1_burstcount),
      .m1_byteenable    (pipeline_bridge_m1_byteenable),
      .m1_chipselect    (pipeline_bridge_m1_chipselect),
      .m1_debugaccess   (pipeline_bridge_m1_debugaccess),
      .m1_endofpacket   (pipeline_bridge_m1_endofpacket),
      .m1_read          (pipeline_bridge_m1_read),
      .m1_readdata      (pipeline_bridge_m1_readdata),
      .m1_readdatavalid (pipeline_bridge_m1_readdatavalid),
      .m1_waitrequest   (pipeline_bridge_m1_waitrequest),
      .m1_write         (pipeline_bridge_m1_write),
      .m1_writedata     (pipeline_bridge_m1_writedata),
      .reset_n          (pipeline_bridge_s1_reset_n),
      .s1_address       (pipeline_bridge_s1_address),
      .s1_arbiterlock   (pipeline_bridge_s1_arbiterlock),
      .s1_arbiterlock2  (pipeline_bridge_s1_arbiterlock2),
      .s1_burstcount    (pipeline_bridge_s1_burstcount),
      .s1_byteenable    (pipeline_bridge_s1_byteenable),
      .s1_chipselect    (pipeline_bridge_s1_chipselect),
      .s1_debugaccess   (pipeline_bridge_s1_debugaccess),
      .s1_endofpacket   (pipeline_bridge_s1_endofpacket),
      .s1_nativeaddress (pipeline_bridge_s1_nativeaddress),
      .s1_read          (pipeline_bridge_s1_read),
      .s1_readdata      (pipeline_bridge_s1_readdata),
      .s1_readdatavalid (pipeline_bridge_s1_readdatavalid),
      .s1_waitrequest   (pipeline_bridge_s1_waitrequest),
      .s1_write         (pipeline_bridge_s1_write),
      .s1_writedata     (pipeline_bridge_s1_writedata)
    );

  push_buttons_s1_arbitrator the_push_buttons_s1
    (
      .clk                                                        (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                  (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_push_buttons_s1           (clock_crossing_bridge_m1_granted_push_buttons_s1),
      .clock_crossing_bridge_m1_latency_counter                   (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                     (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_push_buttons_s1 (clock_crossing_bridge_m1_qualified_request_push_buttons_s1),
      .clock_crossing_bridge_m1_read                              (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_push_buttons_s1   (clock_crossing_bridge_m1_read_data_valid_push_buttons_s1),
      .clock_crossing_bridge_m1_requests_push_buttons_s1          (clock_crossing_bridge_m1_requests_push_buttons_s1),
      .clock_crossing_bridge_m1_write                             (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                         (clock_crossing_bridge_m1_writedata),
      .d1_push_buttons_s1_end_xfer                                (d1_push_buttons_s1_end_xfer),
      .push_buttons_s1_address                                    (push_buttons_s1_address),
      .push_buttons_s1_chipselect                                 (push_buttons_s1_chipselect),
      .push_buttons_s1_irq                                        (push_buttons_s1_irq),
      .push_buttons_s1_irq_from_sa                                (push_buttons_s1_irq_from_sa),
      .push_buttons_s1_readdata                                   (push_buttons_s1_readdata),
      .push_buttons_s1_readdata_from_sa                           (push_buttons_s1_readdata_from_sa),
      .push_buttons_s1_reset_n                                    (push_buttons_s1_reset_n),
      .push_buttons_s1_write_n                                    (push_buttons_s1_write_n),
      .push_buttons_s1_writedata                                  (push_buttons_s1_writedata),
      .reset_n                                                    (slow_clk_reset_n)
    );

  push_buttons the_push_buttons
    (
      .address    (push_buttons_s1_address),
      .chipselect (push_buttons_s1_chipselect),
      .clk        (slow_clk),
      .in_port    (in_port_to_the_push_buttons),
      .irq        (push_buttons_s1_irq),
      .readdata   (push_buttons_s1_readdata),
      .reset_n    (push_buttons_s1_reset_n),
      .write_n    (push_buttons_s1_write_n),
      .writedata  (push_buttons_s1_writedata)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                            (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                      (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_sysid_control_slave           (clock_crossing_bridge_m1_granted_sysid_control_slave),
      .clock_crossing_bridge_m1_latency_counter                       (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                         (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_sysid_control_slave (clock_crossing_bridge_m1_qualified_request_sysid_control_slave),
      .clock_crossing_bridge_m1_read                                  (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_sysid_control_slave   (clock_crossing_bridge_m1_read_data_valid_sysid_control_slave),
      .clock_crossing_bridge_m1_requests_sysid_control_slave          (clock_crossing_bridge_m1_requests_sysid_control_slave),
      .clock_crossing_bridge_m1_write                                 (clock_crossing_bridge_m1_write),
      .d1_sysid_control_slave_end_xfer                                (d1_sysid_control_slave_end_xfer),
      .reset_n                                                        (slow_clk_reset_n),
      .sysid_control_slave_address                                    (sysid_control_slave_address),
      .sysid_control_slave_readdata                                   (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                           (sysid_control_slave_readdata_from_sa),
      .sysid_control_slave_reset_n                                    (sysid_control_slave_reset_n)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .clock    (sysid_control_slave_clock),
      .readdata (sysid_control_slave_readdata),
      .reset_n  (sysid_control_slave_reset_n)
    );

  system_tick_s1_arbitrator the_system_tick_s1
    (
      .clk                                                       (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                 (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_system_tick_s1           (clock_crossing_bridge_m1_granted_system_tick_s1),
      .clock_crossing_bridge_m1_latency_counter                  (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                    (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_system_tick_s1 (clock_crossing_bridge_m1_qualified_request_system_tick_s1),
      .clock_crossing_bridge_m1_read                             (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_system_tick_s1   (clock_crossing_bridge_m1_read_data_valid_system_tick_s1),
      .clock_crossing_bridge_m1_requests_system_tick_s1          (clock_crossing_bridge_m1_requests_system_tick_s1),
      .clock_crossing_bridge_m1_write                            (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                        (clock_crossing_bridge_m1_writedata),
      .d1_system_tick_s1_end_xfer                                (d1_system_tick_s1_end_xfer),
      .reset_n                                                   (slow_clk_reset_n),
      .system_tick_s1_address                                    (system_tick_s1_address),
      .system_tick_s1_chipselect                                 (system_tick_s1_chipselect),
      .system_tick_s1_irq                                        (system_tick_s1_irq),
      .system_tick_s1_irq_from_sa                                (system_tick_s1_irq_from_sa),
      .system_tick_s1_readdata                                   (system_tick_s1_readdata),
      .system_tick_s1_readdata_from_sa                           (system_tick_s1_readdata_from_sa),
      .system_tick_s1_reset_n                                    (system_tick_s1_reset_n),
      .system_tick_s1_write_n                                    (system_tick_s1_write_n),
      .system_tick_s1_writedata                                  (system_tick_s1_writedata)
    );

  system_tick the_system_tick
    (
      .address    (system_tick_s1_address),
      .chipselect (system_tick_s1_chipselect),
      .clk        (slow_clk),
      .irq        (system_tick_s1_irq),
      .readdata   (system_tick_s1_readdata),
      .reset_n    (system_tick_s1_reset_n),
      .write_n    (system_tick_s1_write_n),
      .writedata  (system_tick_s1_writedata)
    );

  touchPanel_irq_n_s1_arbitrator the_touchPanel_irq_n_s1
    (
      .clk                                                            (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                      (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1           (clock_crossing_bridge_m1_granted_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_latency_counter                       (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                         (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1 (clock_crossing_bridge_m1_qualified_request_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_read                                  (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1   (clock_crossing_bridge_m1_read_data_valid_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1          (clock_crossing_bridge_m1_requests_touchPanel_irq_n_s1),
      .clock_crossing_bridge_m1_write                                 (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                             (clock_crossing_bridge_m1_writedata),
      .d1_touchPanel_irq_n_s1_end_xfer                                (d1_touchPanel_irq_n_s1_end_xfer),
      .reset_n                                                        (slow_clk_reset_n),
      .touchPanel_irq_n_s1_address                                    (touchPanel_irq_n_s1_address),
      .touchPanel_irq_n_s1_chipselect                                 (touchPanel_irq_n_s1_chipselect),
      .touchPanel_irq_n_s1_irq                                        (touchPanel_irq_n_s1_irq),
      .touchPanel_irq_n_s1_irq_from_sa                                (touchPanel_irq_n_s1_irq_from_sa),
      .touchPanel_irq_n_s1_readdata                                   (touchPanel_irq_n_s1_readdata),
      .touchPanel_irq_n_s1_readdata_from_sa                           (touchPanel_irq_n_s1_readdata_from_sa),
      .touchPanel_irq_n_s1_reset_n                                    (touchPanel_irq_n_s1_reset_n),
      .touchPanel_irq_n_s1_write_n                                    (touchPanel_irq_n_s1_write_n),
      .touchPanel_irq_n_s1_writedata                                  (touchPanel_irq_n_s1_writedata)
    );

  touchPanel_irq_n the_touchPanel_irq_n
    (
      .address    (touchPanel_irq_n_s1_address),
      .chipselect (touchPanel_irq_n_s1_chipselect),
      .clk        (slow_clk),
      .in_port    (in_port_to_the_touchPanel_irq_n),
      .irq        (touchPanel_irq_n_s1_irq),
      .readdata   (touchPanel_irq_n_s1_readdata),
      .reset_n    (touchPanel_irq_n_s1_reset_n),
      .write_n    (touchPanel_irq_n_s1_write_n),
      .writedata  (touchPanel_irq_n_s1_writedata)
    );

  touchPanel_spi_spi_control_port_arbitrator the_touchPanel_spi_spi_control_port
    (
      .clk                                                                        (slow_clk),
      .clock_crossing_bridge_m1_address_to_slave                                  (clock_crossing_bridge_m1_address_to_slave),
      .clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port           (clock_crossing_bridge_m1_granted_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_latency_counter                                   (clock_crossing_bridge_m1_latency_counter),
      .clock_crossing_bridge_m1_nativeaddress                                     (clock_crossing_bridge_m1_nativeaddress),
      .clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port (clock_crossing_bridge_m1_qualified_request_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_read                                              (clock_crossing_bridge_m1_read),
      .clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port   (clock_crossing_bridge_m1_read_data_valid_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port          (clock_crossing_bridge_m1_requests_touchPanel_spi_spi_control_port),
      .clock_crossing_bridge_m1_write                                             (clock_crossing_bridge_m1_write),
      .clock_crossing_bridge_m1_writedata                                         (clock_crossing_bridge_m1_writedata),
      .d1_touchPanel_spi_spi_control_port_end_xfer                                (d1_touchPanel_spi_spi_control_port_end_xfer),
      .reset_n                                                                    (slow_clk_reset_n),
      .touchPanel_spi_spi_control_port_address                                    (touchPanel_spi_spi_control_port_address),
      .touchPanel_spi_spi_control_port_chipselect                                 (touchPanel_spi_spi_control_port_chipselect),
      .touchPanel_spi_spi_control_port_dataavailable                              (touchPanel_spi_spi_control_port_dataavailable),
      .touchPanel_spi_spi_control_port_dataavailable_from_sa                      (touchPanel_spi_spi_control_port_dataavailable_from_sa),
      .touchPanel_spi_spi_control_port_endofpacket                                (touchPanel_spi_spi_control_port_endofpacket),
      .touchPanel_spi_spi_control_port_endofpacket_from_sa                        (touchPanel_spi_spi_control_port_endofpacket_from_sa),
      .touchPanel_spi_spi_control_port_irq                                        (touchPanel_spi_spi_control_port_irq),
      .touchPanel_spi_spi_control_port_irq_from_sa                                (touchPanel_spi_spi_control_port_irq_from_sa),
      .touchPanel_spi_spi_control_port_read_n                                     (touchPanel_spi_spi_control_port_read_n),
      .touchPanel_spi_spi_control_port_readdata                                   (touchPanel_spi_spi_control_port_readdata),
      .touchPanel_spi_spi_control_port_readdata_from_sa                           (touchPanel_spi_spi_control_port_readdata_from_sa),
      .touchPanel_spi_spi_control_port_readyfordata                               (touchPanel_spi_spi_control_port_readyfordata),
      .touchPanel_spi_spi_control_port_readyfordata_from_sa                       (touchPanel_spi_spi_control_port_readyfordata_from_sa),
      .touchPanel_spi_spi_control_port_reset_n                                    (touchPanel_spi_spi_control_port_reset_n),
      .touchPanel_spi_spi_control_port_write_n                                    (touchPanel_spi_spi_control_port_write_n),
      .touchPanel_spi_spi_control_port_writedata                                  (touchPanel_spi_spi_control_port_writedata)
    );

  touchPanel_spi the_touchPanel_spi
    (
      .MISO          (MISO_to_the_touchPanel_spi),
      .MOSI          (MOSI_from_the_touchPanel_spi),
      .SCLK          (SCLK_from_the_touchPanel_spi),
      .SS_n          (SS_n_from_the_touchPanel_spi),
      .clk           (slow_clk),
      .data_from_cpu (touchPanel_spi_spi_control_port_writedata),
      .data_to_cpu   (touchPanel_spi_spi_control_port_readdata),
      .dataavailable (touchPanel_spi_spi_control_port_dataavailable),
      .endofpacket   (touchPanel_spi_spi_control_port_endofpacket),
      .irq           (touchPanel_spi_spi_control_port_irq),
      .mem_addr      (touchPanel_spi_spi_control_port_address),
      .read_n        (touchPanel_spi_spi_control_port_read_n),
      .readyfordata  (touchPanel_spi_spi_control_port_readyfordata),
      .reset_n       (touchPanel_spi_spi_control_port_reset_n),
      .spi_select    (touchPanel_spi_spi_control_port_chipselect),
      .write_n       (touchPanel_spi_spi_control_port_write_n)
    );

  tristate_bridge_avalon_slave_arbitrator the_tristate_bridge_avalon_slave
    (
      .adsc_n_to_the_ssram                                       (adsc_n_to_the_ssram),
      .bw_n_to_the_ssram                                         (bw_n_to_the_ssram),
      .bwe_n_to_the_ssram                                        (bwe_n_to_the_ssram),
      .chipenable1_n_to_the_ssram                                (chipenable1_n_to_the_ssram),
      .clk                                                       (system_clk),
      .d1_tristate_bridge_avalon_slave_end_xfer                  (d1_tristate_bridge_avalon_slave_end_xfer),
      .flash_s1_wait_counter_eq_0                                (flash_s1_wait_counter_eq_0),
      .flash_ssram_pipeline_bridge_m1_address_to_slave           (flash_ssram_pipeline_bridge_m1_address_to_slave),
      .flash_ssram_pipeline_bridge_m1_burstcount                 (flash_ssram_pipeline_bridge_m1_burstcount),
      .flash_ssram_pipeline_bridge_m1_byteenable                 (flash_ssram_pipeline_bridge_m1_byteenable),
      .flash_ssram_pipeline_bridge_m1_byteenable_flash_s1        (flash_ssram_pipeline_bridge_m1_byteenable_flash_s1),
      .flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1        (flash_ssram_pipeline_bridge_m1_byteenable_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_chipselect                 (flash_ssram_pipeline_bridge_m1_chipselect),
      .flash_ssram_pipeline_bridge_m1_dbs_address                (flash_ssram_pipeline_bridge_m1_dbs_address),
      .flash_ssram_pipeline_bridge_m1_dbs_write_16               (flash_ssram_pipeline_bridge_m1_dbs_write_16),
      .flash_ssram_pipeline_bridge_m1_dbs_write_32               (flash_ssram_pipeline_bridge_m1_dbs_write_32),
      .flash_ssram_pipeline_bridge_m1_granted_flash_s1           (flash_ssram_pipeline_bridge_m1_granted_flash_s1),
      .flash_ssram_pipeline_bridge_m1_granted_ssram_s1           (flash_ssram_pipeline_bridge_m1_granted_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_latency_counter            (flash_ssram_pipeline_bridge_m1_latency_counter),
      .flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1 (flash_ssram_pipeline_bridge_m1_qualified_request_flash_s1),
      .flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1 (flash_ssram_pipeline_bridge_m1_qualified_request_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_read                       (flash_ssram_pipeline_bridge_m1_read),
      .flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1   (flash_ssram_pipeline_bridge_m1_read_data_valid_flash_s1),
      .flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1   (flash_ssram_pipeline_bridge_m1_read_data_valid_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_requests_flash_s1          (flash_ssram_pipeline_bridge_m1_requests_flash_s1),
      .flash_ssram_pipeline_bridge_m1_requests_ssram_s1          (flash_ssram_pipeline_bridge_m1_requests_ssram_s1),
      .flash_ssram_pipeline_bridge_m1_write                      (flash_ssram_pipeline_bridge_m1_write),
      .incoming_tristate_bridge_data                             (incoming_tristate_bridge_data),
      .incoming_tristate_bridge_data_with_Xs_converted_to_0      (incoming_tristate_bridge_data_with_Xs_converted_to_0),
      .outputenable_n_to_the_ssram                               (outputenable_n_to_the_ssram),
      .read_n_to_the_flash                                       (read_n_to_the_flash),
      .reset_n                                                   (system_clk_reset_n),
      .reset_n_to_the_ssram                                      (reset_n_to_the_ssram),
      .select_n_to_the_flash                                     (select_n_to_the_flash),
      .tristate_bridge_address                                   (tristate_bridge_address),
      .tristate_bridge_data                                      (tristate_bridge_data),
      .write_n_to_the_flash                                      (write_n_to_the_flash)
    );

  //reset is asserted asynchronously and deasserted synchronously
  system_reset_system_clk_domain_synch_module system_reset_system_clk_domain_synch
    (
      .clk      (system_clk),
      .data_in  (1'b1),
      .data_out (system_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  system_reset_frame_buffer_phy_clk_out_domain_synch_module system_reset_frame_buffer_phy_clk_out_domain_synch
    (
      .clk      (frame_buffer_phy_clk_out),
      .data_in  (1'b1),
      .data_out (frame_buffer_phy_clk_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  system_reset_slow_clk_domain_synch_module system_reset_slow_clk_domain_synch
    (
      .clk      (slow_clk),
      .data_in  (1'b1),
      .data_out (slow_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  system_reset_video_clk_domain_synch_module system_reset_video_clk_domain_synch
    (
      .clk      (video_clk),
      .data_in  (1'b1),
      .data_out (video_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //ddr_sdram_clock_crossing_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign ddr_sdram_clock_crossing_bridge_m1_endofpacket = 0;

  //flash_ssram_pipeline_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign flash_ssram_pipeline_bridge_m1_endofpacket = 0;

  //sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  assign sysid_control_slave_clock = 0;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_lane0_module (
                            // inputs:
                             data,
                             rdaddress,
                             rdclken,
                             wraddress,
                             wrclock,
                             wren,

                            // outputs:
                             q
                          )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 22: 0] rdaddress;
  input            rdclken;
  input   [ 22: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [8388607: 0];
  wire    [  7: 0] q;
  reg     [ 22: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("flash_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "flash_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 23,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_lane1_module (
                            // inputs:
                             data,
                             rdaddress,
                             rdclken,
                             wraddress,
                             wrclock,
                             wren,

                            // outputs:
                             q
                          )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 22: 0] rdaddress;
  input            rdclken;
  input   [ 22: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [8388607: 0];
  wire    [  7: 0] q;
  reg     [ 22: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("flash_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "flash_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 23,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash (
               // inputs:
                address,
                read_n,
                select_n,
                write_n,

               // outputs:
                data
             )
;

  inout   [ 15: 0] data;
  input   [ 22: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 15: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [ 15: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //flash_lane0, which is an e_ram
  flash_lane0_module flash_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //flash_lane1, which is an e_ram
  flash_lane1_module flash_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? {q_1,
    q_0}: {16{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ssram_lane0_module (
                            // inputs:
                             clk,
                             data,
                             rdaddress,
                             rdclken,
                             reset_n,
                             wraddress,
                             wrclock,
                             wren,

                            // outputs:
                             q
                          )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 17: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ssram_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ssram_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ssram_lane1_module (
                            // inputs:
                             clk,
                             data,
                             rdaddress,
                             rdclken,
                             reset_n,
                             wraddress,
                             wrclock,
                             wren,

                            // outputs:
                             q
                          )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 17: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ssram_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ssram_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ssram_lane2_module (
                            // inputs:
                             clk,
                             data,
                             rdaddress,
                             rdclken,
                             reset_n,
                             wraddress,
                             wrclock,
                             wren,

                            // outputs:
                             q
                          )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 17: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ssram_lane2.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ssram_lane2.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ssram_lane3_module (
                            // inputs:
                             clk,
                             data,
                             rdaddress,
                             rdclken,
                             reset_n,
                             wraddress,
                             wrclock,
                             wren,

                            // outputs:
                             q
                          )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 17: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 17: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 17: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [262143: 0];
  wire    [  7: 0] q;
  reg     [ 17: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ssram_lane3.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ssram_lane3.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 18,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ssram (
               // inputs:
                address,
                adsc_n,
                bw_n,
                bwe_n,
                chipenable1_n,
                clk,
                outputenable_n,
                reset_n,

               // outputs:
                data
             )
;

  inout   [ 31: 0] data;
  input   [ 17: 0] address;
  input            adsc_n;
  input   [  3: 0] bw_n;
  input            bwe_n;
  input            chipenable1_n;
  input            clk;
  input            outputenable_n;
  input            reset_n;

  wire    [ 31: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [  7: 0] data_2;
  wire    [  7: 0] data_3;
  wire    [ 31: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  wire    [  7: 0] q_2;
  wire    [  7: 0] q_3;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ssram_lane0, which is an e_ram
  ssram_lane0_module ssram_lane0
    (
      .clk       (clk),
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[0])
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ssram_lane1, which is an e_ram
  ssram_lane1_module ssram_lane1
    (
      .clk       (clk),
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[1])
    );

  assign data_2 = logic_vector_gasket[23 : 16];
  //ssram_lane2, which is an e_ram
  ssram_lane2_module ssram_lane2
    (
      .clk       (clk),
      .data      (data_2),
      .q         (q_2),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[2])
    );

  assign data_3 = logic_vector_gasket[31 : 24];
  //ssram_lane3, which is an e_ram
  ssram_lane3_module ssram_lane3
    (
      .clk       (clk),
      .data      (data_3),
      .q         (q_3),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[3])
    );

  assign data = (~chipenable1_n & ~outputenable_n)? {q_3,
    q_2,
    q_1,
    q_0}: {32{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "d:/altera/12.1/quartus/eda/sim_lib/altera_mf.v"
`include "d:/altera/12.1/quartus/eda/sim_lib/220model.v"
`include "d:/altera/12.1/quartus/eda/sim_lib/sgate.v"
`include "accelerator_mandelbrot_hw_draw_int_mandelbrot.v"
`include "accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance.v"
`include "dummy_master/dummy_master.v"
`include "dummy_master_inst.v"
`include "lcd_pixel_converter.vo"
`include "lcd_video_sequencer.vo"
`include "descriptor_memory.v"
`include "sysid.v"
`include "colour_lookup_table.v"
`include "pio_id_eeprom_scl.v"
`include "push_buttons.v"
`include "jtag_uart.v"
`include "lcd_ta_formatter_to_fifo.v"
`include "pipeline_bridge.v"
`include "pio_id_eeprom_dat.v"
`include "lcd_ta_fifo_to_sequencer.v"
`include "lcd_ta_fifo_to_sequencer_fifo.v"
`include "cpu_test_bench.v"
`include "cpu_mult_cell.v"
`include "cpu_oci_test_bench.v"
`include "cpu_jtag_debug_module_tck.v"
`include "cpu_jtag_debug_module_sysclk.v"
`include "cpu_jtag_debug_module_wrapper.v"
`include "cpu.v"
`include "lcd_data_format_adapter.v"
`include "lcd_data_format_adapter_state_ram.v"
`include "lcd_data_format_adapter_data_ram.v"
`include "lcd_on_chip_memory_fifo.v"
`include "lcd_sgdma.v"
`include "clock_crossing_bridge.v"
`include "lcd_i2c_dat.v"
`include "lcd_i2c_scl.v"
`include "touchPanel_spi.v"
`include "system_tick.v"
`include "lcd_i2c_cs.v"
`include "frame_buffer_pipeline_bridge.v"
`include "touchPanel_irq_n.v"
`include "lcd_data_format_adapter_1.v"
`include "flash_ssram_pipeline_bridge.v"
`include "ddr_sdram_clock_crossing_bridge.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire             DEN_from_the_lcd_video_sequencer;
  wire             HD_from_the_lcd_video_sequencer;
  wire             MISO_to_the_touchPanel_spi;
  wire             MOSI_from_the_touchPanel_spi;
  wire    [  7: 0] RGB_OUT_from_the_lcd_video_sequencer;
  wire             SCLK_from_the_touchPanel_spi;
  wire             SS_n_from_the_touchPanel_spi;
  wire             VD_from_the_lcd_video_sequencer;
  wire    [ 31: 0] accelerator_mandelbrot_hw_draw_int_mandelbrot_managed_instance_dummy_slave_readdata_from_sa;
  wire             adsc_n_to_the_ssram;
  wire             bidir_port_to_and_from_the_lcd_i2c_dat;
  wire             bidir_port_to_and_from_the_pio_id_eeprom_dat;
  wire    [  3: 0] bw_n_to_the_ssram;
  wire             bwe_n_to_the_ssram;
  wire             chipenable1_n_to_the_ssram;
  wire             clk;
  wire             ddr_sdram_clock_crossing_bridge_m1_endofpacket;
  wire    [ 22: 0] ddr_sdram_clock_crossing_bridge_m1_nativeaddress;
  reg              ext_clk_one;
  wire             flash_ssram_pipeline_bridge_m1_debugaccess;
  wire             flash_ssram_pipeline_bridge_m1_endofpacket;
  wire             frame_buffer_aux_full_rate_clk_out;
  wire             frame_buffer_aux_half_rate_clk_out;
  wire             frame_buffer_phy_clk_out;
  wire             frame_buffer_pipeline_bridge_m1_debugaccess;
  wire             global_reset_n_to_the_frame_buffer;
  wire    [  3: 0] in_port_to_the_push_buttons;
  wire             in_port_to_the_touchPanel_irq_n;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             local_init_done_from_the_frame_buffer;
  wire             local_refresh_ack_from_the_frame_buffer;
  wire             local_wdata_req_from_the_frame_buffer;
  wire    [ 12: 0] mem_addr_from_the_frame_buffer;
  wire    [  1: 0] mem_ba_from_the_frame_buffer;
  wire             mem_cas_n_from_the_frame_buffer;
  wire             mem_cke_from_the_frame_buffer;
  wire             mem_clk_n_to_and_from_the_frame_buffer;
  wire             mem_clk_to_and_from_the_frame_buffer;
  wire             mem_cs_n_from_the_frame_buffer;
  wire    [  1: 0] mem_dm_from_the_frame_buffer;
  wire    [ 15: 0] mem_dq_to_and_from_the_frame_buffer;
  wire    [  1: 0] mem_dqs_to_and_from_the_frame_buffer;
  wire             mem_ras_n_from_the_frame_buffer;
  wire             mem_we_n_from_the_frame_buffer;
  wire             out_port_from_the_lcd_i2c_cs;
  wire             out_port_from_the_lcd_i2c_scl;
  wire             out_port_from_the_pio_id_eeprom_scl;
  wire             outputenable_n_to_the_ssram;
  wire             pipeline_bridge_s1_endofpacket_from_sa;
  wire             read_n_to_the_flash;
  reg              reset_n;
  wire             reset_n_to_the_ssram;
  wire             reset_phy_clk_n_from_the_frame_buffer;
  wire             select_n_to_the_flash;
  reg              slow_clk;
  wire             sysid_control_slave_clock;
  reg              system_clk;
  wire             touchPanel_spi_spi_control_port_dataavailable_from_sa;
  wire             touchPanel_spi_spi_control_port_readyfordata_from_sa;
  wire    [ 23: 0] tristate_bridge_address;
  wire    [ 31: 0] tristate_bridge_data;
  reg              video_clk;
  wire             write_n_to_the_flash;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  system DUT
    (
      .DEN_from_the_lcd_video_sequencer             (DEN_from_the_lcd_video_sequencer),
      .HD_from_the_lcd_video_sequencer              (HD_from_the_lcd_video_sequencer),
      .MISO_to_the_touchPanel_spi                   (MISO_to_the_touchPanel_spi),
      .MOSI_from_the_touchPanel_spi                 (MOSI_from_the_touchPanel_spi),
      .RGB_OUT_from_the_lcd_video_sequencer         (RGB_OUT_from_the_lcd_video_sequencer),
      .SCLK_from_the_touchPanel_spi                 (SCLK_from_the_touchPanel_spi),
      .SS_n_from_the_touchPanel_spi                 (SS_n_from_the_touchPanel_spi),
      .VD_from_the_lcd_video_sequencer              (VD_from_the_lcd_video_sequencer),
      .adsc_n_to_the_ssram                          (adsc_n_to_the_ssram),
      .bidir_port_to_and_from_the_lcd_i2c_dat       (bidir_port_to_and_from_the_lcd_i2c_dat),
      .bidir_port_to_and_from_the_pio_id_eeprom_dat (bidir_port_to_and_from_the_pio_id_eeprom_dat),
      .bw_n_to_the_ssram                            (bw_n_to_the_ssram),
      .bwe_n_to_the_ssram                           (bwe_n_to_the_ssram),
      .chipenable1_n_to_the_ssram                   (chipenable1_n_to_the_ssram),
      .ext_clk_one                                  (ext_clk_one),
      .frame_buffer_aux_full_rate_clk_out           (frame_buffer_aux_full_rate_clk_out),
      .frame_buffer_aux_half_rate_clk_out           (frame_buffer_aux_half_rate_clk_out),
      .frame_buffer_phy_clk_out                     (frame_buffer_phy_clk_out),
      .global_reset_n_to_the_frame_buffer           (global_reset_n_to_the_frame_buffer),
      .in_port_to_the_push_buttons                  (in_port_to_the_push_buttons),
      .in_port_to_the_touchPanel_irq_n              (in_port_to_the_touchPanel_irq_n),
      .local_init_done_from_the_frame_buffer        (local_init_done_from_the_frame_buffer),
      .local_refresh_ack_from_the_frame_buffer      (local_refresh_ack_from_the_frame_buffer),
      .local_wdata_req_from_the_frame_buffer        (local_wdata_req_from_the_frame_buffer),
      .mem_addr_from_the_frame_buffer               (mem_addr_from_the_frame_buffer),
      .mem_ba_from_the_frame_buffer                 (mem_ba_from_the_frame_buffer),
      .mem_cas_n_from_the_frame_buffer              (mem_cas_n_from_the_frame_buffer),
      .mem_cke_from_the_frame_buffer                (mem_cke_from_the_frame_buffer),
      .mem_clk_n_to_and_from_the_frame_buffer       (mem_clk_n_to_and_from_the_frame_buffer),
      .mem_clk_to_and_from_the_frame_buffer         (mem_clk_to_and_from_the_frame_buffer),
      .mem_cs_n_from_the_frame_buffer               (mem_cs_n_from_the_frame_buffer),
      .mem_dm_from_the_frame_buffer                 (mem_dm_from_the_frame_buffer),
      .mem_dq_to_and_from_the_frame_buffer          (mem_dq_to_and_from_the_frame_buffer),
      .mem_dqs_to_and_from_the_frame_buffer         (mem_dqs_to_and_from_the_frame_buffer),
      .mem_ras_n_from_the_frame_buffer              (mem_ras_n_from_the_frame_buffer),
      .mem_we_n_from_the_frame_buffer               (mem_we_n_from_the_frame_buffer),
      .out_port_from_the_lcd_i2c_cs                 (out_port_from_the_lcd_i2c_cs),
      .out_port_from_the_lcd_i2c_scl                (out_port_from_the_lcd_i2c_scl),
      .out_port_from_the_pio_id_eeprom_scl          (out_port_from_the_pio_id_eeprom_scl),
      .outputenable_n_to_the_ssram                  (outputenable_n_to_the_ssram),
      .read_n_to_the_flash                          (read_n_to_the_flash),
      .reset_n                                      (reset_n),
      .reset_n_to_the_ssram                         (reset_n_to_the_ssram),
      .reset_phy_clk_n_from_the_frame_buffer        (reset_phy_clk_n_from_the_frame_buffer),
      .select_n_to_the_flash                        (select_n_to_the_flash),
      .slow_clk                                     (slow_clk),
      .system_clk                                   (system_clk),
      .tristate_bridge_address                      (tristate_bridge_address),
      .tristate_bridge_data                         (tristate_bridge_data),
      .video_clk                                    (video_clk),
      .write_n_to_the_flash                         (write_n_to_the_flash)
    );

  flash the_flash
    (
      .address  (tristate_bridge_address[23 : 1]),
      .data     (tristate_bridge_data),
      .read_n   (read_n_to_the_flash),
      .select_n (select_n_to_the_flash),
      .write_n  (write_n_to_the_flash)
    );

  //default value specified in MODULE push_buttons ptf port section
  assign in_port_to_the_push_buttons = 15;

  ssram the_ssram
    (
      .address        (tristate_bridge_address[19 : 2]),
      .adsc_n         (adsc_n_to_the_ssram),
      .bw_n           (bw_n_to_the_ssram),
      .bwe_n          (bwe_n_to_the_ssram),
      .chipenable1_n  (chipenable1_n_to_the_ssram),
      .clk            (system_clk),
      .data           (tristate_bridge_data),
      .outputenable_n (outputenable_n_to_the_ssram),
      .reset_n        (reset_n_to_the_ssram)
    );

  initial
    ext_clk_one = 1'b0;
  always
    #10 ext_clk_one <= ~ext_clk_one;
  
  initial 
    begin
      reset_n <= 0;
      #200 reset_n <= 1;
    end
  initial
    slow_clk = 1'b0;
  always
    #10 slow_clk <= ~slow_clk;
  
  initial
    system_clk = 1'b0;
  always
    #5 system_clk <= ~system_clk;
  
  initial
    video_clk = 1'b0;
  always
    #5 video_clk <= ~video_clk;
  

endmodule


//synthesis translate_on